

module Stat_2000_304
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1922,
  n1924,
  n1926,
  n1925,
  n1957,
  n1952,
  n1943,
  n1951,
  n1946,
  n1944,
  n1955,
  n1948,
  n1971,
  n1966,
  n1967,
  n1969,
  n1974,
  n2023,
  n2020,
  n2028,
  n2027,
  n2021,
  n2025,
  n2032,
  n2019,
  n2030,
  n2018,
  n2031,
  n2022,
  n2024,
  n2026,
  n2029
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n1922;output n1924;output n1926;output n1925;output n1957;output n1952;output n1943;output n1951;output n1946;output n1944;output n1955;output n1948;output n1971;output n1966;output n1967;output n1969;output n1974;output n2023;output n2020;output n2028;output n2027;output n2021;output n2025;output n2032;output n2019;output n2030;output n2018;output n2031;output n2022;output n2024;output n2026;output n2029;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1923;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1945;wire n1947;wire n1949;wire n1950;wire n1953;wire n1954;wire n1956;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1968;wire n1970;wire n1972;wire n1973;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;

  buf
  g0
  (
    n47,
    n6
  );


  buf
  g1
  (
    n44,
    n3
  );


  not
  g2
  (
    n40,
    n5
  );


  not
  g3
  (
    n37,
    n2
  );


  buf
  g4
  (
    n43,
    n6
  );


  buf
  g5
  (
    n42,
    n4
  );


  not
  g6
  (
    n41,
    n1
  );


  buf
  g7
  (
    n39,
    n4
  );


  not
  g8
  (
    n36,
    n2
  );


  buf
  g9
  (
    n46,
    n3
  );


  not
  g10
  (
    n33,
    n5
  );


  buf
  g11
  (
    n38,
    n6
  );


  buf
  g12
  (
    n45,
    n5
  );


  buf
  g13
  (
    n35,
    n5
  );


  not
  g14
  (
    n48,
    n1
  );


  buf
  g15
  (
    n53,
    n2
  );


  not
  g16
  (
    n55,
    n2
  );


  not
  g17
  (
    n50,
    n1
  );


  buf
  g18
  (
    n34,
    n3
  );


  buf
  g19
  (
    n52,
    n3
  );


  not
  g20
  (
    n54,
    n4
  );


  not
  g21
  (
    n51,
    n4
  );


  not
  g22
  (
    n49,
    n1
  );


  buf
  g23
  (
    n111,
    n43
  );


  not
  g24
  (
    n88,
    n34
  );


  not
  g25
  (
    n114,
    n36
  );


  buf
  g26
  (
    n81,
    n42
  );


  buf
  g27
  (
    n79,
    n34
  );


  not
  g28
  (
    n65,
    n44
  );


  buf
  g29
  (
    KeyWire_0_2,
    n34
  );


  buf
  g30
  (
    n73,
    n42
  );


  buf
  g31
  (
    n101,
    n48
  );


  buf
  g32
  (
    n69,
    n38
  );


  buf
  g33
  (
    n118,
    n46
  );


  not
  g34
  (
    n91,
    n34
  );


  not
  g35
  (
    n92,
    n33
  );


  not
  g36
  (
    n67,
    n44
  );


  buf
  g37
  (
    n120,
    n48
  );


  not
  g38
  (
    n62,
    n45
  );


  not
  g39
  (
    n76,
    n47
  );


  not
  g40
  (
    n103,
    n39
  );


  not
  g41
  (
    n78,
    n42
  );


  buf
  g42
  (
    n97,
    n33
  );


  not
  g43
  (
    n94,
    n50
  );


  buf
  g44
  (
    n61,
    n35
  );


  buf
  g45
  (
    n102,
    n50
  );


  buf
  g46
  (
    n63,
    n47
  );


  not
  g47
  (
    n66,
    n43
  );


  not
  g48
  (
    n56,
    n49
  );


  buf
  g49
  (
    n83,
    n35
  );


  buf
  g50
  (
    n90,
    n41
  );


  not
  g51
  (
    n89,
    n44
  );


  buf
  g52
  (
    n116,
    n43
  );


  buf
  g53
  (
    n119,
    n37
  );


  not
  g54
  (
    n98,
    n38
  );


  buf
  g55
  (
    n68,
    n38
  );


  buf
  g56
  (
    n99,
    n44
  );


  buf
  g57
  (
    n110,
    n37
  );


  buf
  g58
  (
    n100,
    n42
  );


  buf
  g59
  (
    n95,
    n46
  );


  not
  g60
  (
    n106,
    n47
  );


  not
  g61
  (
    n72,
    n40
  );


  not
  g62
  (
    n82,
    n46
  );


  buf
  g63
  (
    n96,
    n48
  );


  buf
  g64
  (
    n87,
    n49
  );


  buf
  g65
  (
    n70,
    n48
  );


  not
  g66
  (
    n74,
    n45
  );


  not
  g67
  (
    n60,
    n45
  );


  not
  g68
  (
    n121,
    n41
  );


  buf
  g69
  (
    n57,
    n39
  );


  buf
  g70
  (
    n80,
    n36
  );


  buf
  g71
  (
    n104,
    n33
  );


  buf
  g72
  (
    n108,
    n49
  );


  not
  g73
  (
    n109,
    n46
  );


  buf
  g74
  (
    n112,
    n40
  );


  buf
  g75
  (
    n75,
    n39
  );


  buf
  g76
  (
    n64,
    n33
  );


  buf
  g77
  (
    n58,
    n43
  );


  buf
  g78
  (
    n84,
    n47
  );


  not
  g79
  (
    n105,
    n36
  );


  buf
  g80
  (
    n77,
    n50
  );


  buf
  g81
  (
    n113,
    n40
  );


  not
  g82
  (
    n59,
    n38
  );


  not
  g83
  (
    n86,
    n49
  );


  nor
  g84
  (
    n85,
    n39,
    n37
  );


  xnor
  g85
  (
    n115,
    n35,
    n36
  );


  and
  g86
  (
    n93,
    n37,
    n41
  );


  or
  g87
  (
    n117,
    n41,
    n45
  );


  or
  g88
  (
    n107,
    n35,
    n40
  );


  nor
  g89
  (
    n123,
    n67,
    n63,
    n74,
    n71
  );


  and
  g90
  (
    n127,
    n73,
    n65,
    n61,
    n59
  );


  xnor
  g91
  (
    n124,
    n82,
    n64,
    n86,
    n75
  );


  xnor
  g92
  (
    n126,
    n79,
    n77,
    n56,
    n78
  );


  or
  g93
  (
    n122,
    n87,
    n76,
    n62,
    n69
  );


  xor
  g94
  (
    n125,
    n68,
    n70,
    n58,
    n72
  );


  nand
  g95
  (
    n128,
    n83,
    n85,
    n57,
    n81
  );


  xor
  g96
  (
    n129,
    n60,
    n66,
    n80,
    n84
  );


  not
  g97
  (
    n131,
    n127
  );


  buf
  g98
  (
    n135,
    n125
  );


  not
  g99
  (
    n143,
    n127
  );


  buf
  g100
  (
    n142,
    n128
  );


  not
  g101
  (
    n140,
    n129
  );


  not
  g102
  (
    n134,
    n127
  );


  not
  g103
  (
    n132,
    n127
  );


  not
  g104
  (
    n137,
    n128
  );


  not
  g105
  (
    n130,
    n123
  );


  not
  g106
  (
    n144,
    n128
  );


  not
  g107
  (
    n145,
    n122
  );


  not
  g108
  (
    n136,
    n129
  );


  buf
  g109
  (
    n133,
    n124
  );


  not
  g110
  (
    n141,
    n126
  );


  buf
  g111
  (
    n138,
    n126
  );


  not
  g112
  (
    n139,
    n128
  );


  buf
  g113
  (
    n183,
    n144
  );


  buf
  g114
  (
    n174,
    n134
  );


  buf
  g115
  (
    n156,
    n132
  );


  buf
  g116
  (
    n152,
    n139
  );


  not
  g117
  (
    n168,
    n141
  );


  buf
  g118
  (
    n181,
    n139
  );


  buf
  g119
  (
    n177,
    n145
  );


  not
  g120
  (
    n150,
    n52
  );


  not
  g121
  (
    n188,
    n137
  );


  not
  g122
  (
    n172,
    n138
  );


  not
  g123
  (
    n164,
    n54
  );


  buf
  g124
  (
    n175,
    n53
  );


  buf
  g125
  (
    n173,
    n137
  );


  not
  g126
  (
    n170,
    n138
  );


  buf
  g127
  (
    n184,
    n133
  );


  buf
  g128
  (
    n193,
    n141
  );


  not
  g129
  (
    n179,
    n136
  );


  buf
  g130
  (
    n182,
    n138
  );


  buf
  g131
  (
    n148,
    n142
  );


  not
  g132
  (
    n176,
    n144
  );


  not
  g133
  (
    n158,
    n143
  );


  not
  g134
  (
    n166,
    n131
  );


  buf
  g135
  (
    n165,
    n53
  );


  not
  g136
  (
    n160,
    n145
  );


  not
  g137
  (
    n147,
    n52
  );


  buf
  g138
  (
    KeyWire_0_15,
    n52
  );


  not
  g139
  (
    n169,
    n141
  );


  not
  g140
  (
    n149,
    n50
  );


  not
  g141
  (
    n159,
    n143
  );


  buf
  g142
  (
    n171,
    n51
  );


  not
  g143
  (
    n155,
    n145
  );


  buf
  g144
  (
    n154,
    n139
  );


  buf
  g145
  (
    n151,
    n145
  );


  buf
  g146
  (
    n161,
    n132
  );


  buf
  g147
  (
    n162,
    n143
  );


  not
  g148
  (
    n146,
    n144
  );


  not
  g149
  (
    n190,
    n141
  );


  not
  g150
  (
    n178,
    n143
  );


  not
  g151
  (
    n185,
    n134
  );


  not
  g152
  (
    n157,
    n144
  );


  not
  g153
  (
    n167,
    n52
  );


  and
  g154
  (
    n187,
    n131,
    n142,
    n140
  );


  nand
  g155
  (
    n180,
    n53,
    n142,
    n138
  );


  nor
  g156
  (
    n153,
    n139,
    n140,
    n137
  );


  nand
  g157
  (
    n186,
    n140,
    n54,
    n51
  );


  nand
  g158
  (
    n189,
    n135,
    n142,
    n51
  );


  xor
  g159
  (
    n163,
    n135,
    n53,
    n51
  );


  xor
  g160
  (
    n191,
    n133,
    n136,
    n130,
    n140
  );


  buf
  g161
  (
    n274,
    n166
  );


  not
  g162
  (
    n203,
    n159
  );


  not
  g163
  (
    n240,
    n171
  );


  buf
  g164
  (
    n358,
    n96
  );


  buf
  g165
  (
    n241,
    n178
  );


  buf
  g166
  (
    n195,
    n178
  );


  buf
  g167
  (
    n355,
    n146
  );


  not
  g168
  (
    n303,
    n107
  );


  not
  g169
  (
    n283,
    n106
  );


  not
  g170
  (
    n311,
    n97
  );


  buf
  g171
  (
    n265,
    n165
  );


  buf
  g172
  (
    n337,
    n183
  );


  buf
  g173
  (
    n262,
    n182
  );


  not
  g174
  (
    n305,
    n175
  );


  buf
  g175
  (
    n286,
    n158
  );


  not
  g176
  (
    n257,
    n186
  );


  buf
  g177
  (
    n304,
    n181
  );


  not
  g178
  (
    n260,
    n108
  );


  buf
  g179
  (
    n196,
    n114
  );


  not
  g180
  (
    n295,
    n156
  );


  buf
  g181
  (
    n251,
    n157
  );


  buf
  g182
  (
    n360,
    n105
  );


  not
  g183
  (
    n214,
    n164
  );


  not
  g184
  (
    n200,
    n161
  );


  not
  g185
  (
    n339,
    n117
  );


  not
  g186
  (
    n309,
    n176
  );


  buf
  g187
  (
    KeyWire_0_13,
    n95
  );


  buf
  g188
  (
    n207,
    n104
  );


  not
  g189
  (
    n289,
    n170
  );


  buf
  g190
  (
    n365,
    n108
  );


  not
  g191
  (
    n362,
    n147
  );


  not
  g192
  (
    n316,
    n180
  );


  not
  g193
  (
    n243,
    n155
  );


  buf
  g194
  (
    n220,
    n114
  );


  not
  g195
  (
    n300,
    n188
  );


  not
  g196
  (
    n315,
    n154
  );


  not
  g197
  (
    n352,
    n174
  );


  not
  g198
  (
    n204,
    n181
  );


  not
  g199
  (
    n279,
    n182
  );


  not
  g200
  (
    n273,
    n110
  );


  buf
  g201
  (
    n211,
    n91
  );


  buf
  g202
  (
    n278,
    n160
  );


  not
  g203
  (
    n198,
    n112
  );


  buf
  g204
  (
    n230,
    n167
  );


  not
  g205
  (
    n223,
    n172
  );


  buf
  g206
  (
    n197,
    n157
  );


  buf
  g207
  (
    n314,
    n176
  );


  not
  g208
  (
    n349,
    n148
  );


  buf
  g209
  (
    n326,
    n119
  );


  not
  g210
  (
    n194,
    n170
  );


  not
  g211
  (
    n208,
    n177
  );


  buf
  g212
  (
    n340,
    n116
  );


  not
  g213
  (
    n224,
    n111
  );


  buf
  g214
  (
    n282,
    n179
  );


  not
  g215
  (
    n359,
    n165
  );


  buf
  g216
  (
    n338,
    n166
  );


  buf
  g217
  (
    n357,
    n167
  );


  buf
  g218
  (
    n336,
    n107
  );


  not
  g219
  (
    n284,
    n159
  );


  not
  g220
  (
    n341,
    n162
  );


  not
  g221
  (
    n344,
    n173
  );


  not
  g222
  (
    n330,
    n177
  );


  not
  g223
  (
    n333,
    n168
  );


  not
  g224
  (
    n256,
    n110
  );


  not
  g225
  (
    n285,
    n163
  );


  not
  g226
  (
    n346,
    n174
  );


  not
  g227
  (
    n364,
    n158
  );


  not
  g228
  (
    n293,
    n188
  );


  buf
  g229
  (
    n281,
    n162
  );


  buf
  g230
  (
    n345,
    n104
  );


  buf
  g231
  (
    n332,
    n189
  );


  not
  g232
  (
    n235,
    n119
  );


  not
  g233
  (
    n202,
    n188
  );


  buf
  g234
  (
    n328,
    n147
  );


  buf
  g235
  (
    n237,
    n172
  );


  not
  g236
  (
    n266,
    n55
  );


  not
  g237
  (
    n350,
    n184
  );


  not
  g238
  (
    n353,
    n180
  );


  not
  g239
  (
    n347,
    n104
  );


  buf
  g240
  (
    n297,
    n90
  );


  not
  g241
  (
    n210,
    n146
  );


  buf
  g242
  (
    n298,
    n168
  );


  buf
  g243
  (
    n267,
    n176
  );


  not
  g244
  (
    n218,
    n180
  );


  buf
  g245
  (
    n215,
    n114
  );


  buf
  g246
  (
    n319,
    n187
  );


  buf
  g247
  (
    n250,
    n148
  );


  not
  g248
  (
    n205,
    n103
  );


  buf
  g249
  (
    n331,
    n157
  );


  buf
  g250
  (
    n228,
    n156
  );


  not
  g251
  (
    n369,
    n160
  );


  not
  g252
  (
    n272,
    n165
  );


  not
  g253
  (
    n342,
    n175
  );


  buf
  g254
  (
    n264,
    n110
  );


  not
  g255
  (
    KeyWire_0_9,
    n150
  );


  buf
  g256
  (
    n247,
    n112
  );


  not
  g257
  (
    n233,
    n101
  );


  not
  g258
  (
    n252,
    n54
  );


  not
  g259
  (
    n294,
    n113
  );


  buf
  g260
  (
    n348,
    n189
  );


  not
  g261
  (
    n356,
    n165
  );


  buf
  g262
  (
    KeyWire_0_4,
    n156
  );


  buf
  g263
  (
    n288,
    n155
  );


  not
  g264
  (
    n307,
    n103
  );


  buf
  g265
  (
    n317,
    n148
  );


  buf
  g266
  (
    n335,
    n153
  );


  buf
  g267
  (
    n361,
    n164
  );


  not
  g268
  (
    n292,
    n185
  );


  buf
  g269
  (
    n322,
    n163
  );


  buf
  g270
  (
    n299,
    n187
  );


  not
  g271
  (
    n229,
    n176
  );


  buf
  g272
  (
    n287,
    n107
  );


  not
  g273
  (
    n258,
    n113
  );


  buf
  g274
  (
    n259,
    n173
  );


  not
  g275
  (
    n222,
    n116
  );


  buf
  g276
  (
    n306,
    n115
  );


  buf
  g277
  (
    n323,
    n98
  );


  buf
  g278
  (
    n343,
    n107
  );


  buf
  g279
  (
    n363,
    n166
  );


  not
  g280
  (
    n367,
    n105
  );


  not
  g281
  (
    n231,
    n173
  );


  buf
  g282
  (
    n366,
    n189
  );


  buf
  g283
  (
    n368,
    n93
  );


  buf
  g284
  (
    n321,
    n113
  );


  not
  g285
  (
    n213,
    n169
  );


  buf
  g286
  (
    n291,
    n114
  );


  buf
  g287
  (
    n324,
    n172
  );


  buf
  g288
  (
    n253,
    n112
  );


  buf
  g289
  (
    n312,
    n151
  );


  buf
  g290
  (
    n270,
    n161
  );


  not
  g291
  (
    n354,
    n105
  );


  buf
  g292
  (
    n245,
    n186
  );


  buf
  g293
  (
    n234,
    n111
  );


  not
  g294
  (
    n244,
    n166
  );


  not
  g295
  (
    n329,
    n89
  );


  buf
  g296
  (
    n302,
    n168
  );


  not
  g297
  (
    n301,
    n186
  );


  buf
  g298
  (
    n227,
    n167
  );


  not
  g299
  (
    n238,
    n115
  );


  buf
  g300
  (
    n296,
    n161
  );


  buf
  g301
  (
    n232,
    n187
  );


  not
  g302
  (
    n313,
    n161
  );


  buf
  g303
  (
    n248,
    n169
  );


  buf
  g304
  (
    n217,
    n149
  );


  buf
  g305
  (
    n255,
    n109
  );


  buf
  g306
  (
    n320,
    n168
  );


  not
  g307
  (
    n219,
    n181
  );


  not
  g308
  (
    n199,
    n159
  );


  and
  g309
  (
    n308,
    n99,
    n164
  );


  xor
  g310
  (
    n216,
    n151,
    n171,
    n184,
    n162
  );


  xor
  g311
  (
    n225,
    n115,
    n160,
    n180,
    n164
  );


  and
  g312
  (
    n246,
    n149,
    n185,
    n188,
    n150
  );


  xnor
  g313
  (
    n290,
    n117,
    n109,
    n186,
    n155
  );


  nand
  g314
  (
    n254,
    n181,
    n117,
    n92,
    n153
  );


  nor
  g315
  (
    n327,
    n106,
    n116,
    n148,
    n94
  );


  nor
  g316
  (
    n271,
    n151,
    n106,
    n174,
    n179
  );


  or
  g317
  (
    n242,
    n175,
    n88,
    n169,
    n171
  );


  and
  g318
  (
    n236,
    n102,
    n147,
    n109,
    n146
  );


  xor
  g319
  (
    n268,
    n183,
    n118,
    n170,
    n154
  );


  xnor
  g320
  (
    n310,
    n105,
    n178,
    n171,
    n153
  );


  xor
  g321
  (
    n269,
    n163,
    n155,
    n184,
    n113
  );


  nor
  g322
  (
    n275,
    n173,
    n104,
    n158,
    n149
  );


  xnor
  g323
  (
    n318,
    n177,
    n115,
    n182,
    n175
  );


  xor
  g324
  (
    n261,
    n154,
    n185,
    n118
  );


  or
  g325
  (
    n239,
    n158,
    n152,
    n149,
    n178
  );


  xnor
  g326
  (
    n351,
    n159,
    n151,
    n111,
    n187
  );


  and
  g327
  (
    n280,
    n170,
    n189,
    n153,
    n54
  );


  nand
  g328
  (
    n209,
    n116,
    n117,
    n150,
    n152
  );


  nand
  g329
  (
    n263,
    n179,
    n169,
    n146,
    n109
  );


  xnor
  g330
  (
    n226,
    n152,
    n110,
    n111,
    n167
  );


  nand
  g331
  (
    n325,
    n154,
    n182,
    n184,
    n112
  );


  xnor
  g332
  (
    n206,
    n163,
    n162,
    n100,
    n108
  );


  nor
  g333
  (
    n249,
    n185,
    n106,
    n152,
    n177
  );


  xnor
  g334
  (
    n334,
    n172,
    n160,
    n118,
    n174
  );


  nor
  g335
  (
    n221,
    n150,
    n108,
    n157,
    n179
  );


  xor
  g336
  (
    n201,
    n156,
    n147,
    n183
  );


  buf
  g337
  (
    n624,
    n287
  );


  not
  g338
  (
    n713,
    n292
  );


  not
  g339
  (
    n748,
    n205
  );


  buf
  g340
  (
    n950,
    n267
  );


  not
  g341
  (
    n591,
    n198
  );


  not
  g342
  (
    n452,
    n214
  );


  buf
  g343
  (
    n426,
    n196
  );


  buf
  g344
  (
    n566,
    n327
  );


  buf
  g345
  (
    n750,
    n317
  );


  buf
  g346
  (
    n880,
    n319
  );


  buf
  g347
  (
    n541,
    n342
  );


  not
  g348
  (
    n416,
    n257
  );


  buf
  g349
  (
    n1005,
    n339
  );


  buf
  g350
  (
    n484,
    n333
  );


  buf
  g351
  (
    n840,
    n200
  );


  not
  g352
  (
    n617,
    n337
  );


  not
  g353
  (
    n593,
    n319
  );


  not
  g354
  (
    n638,
    n328
  );


  buf
  g355
  (
    n723,
    n250
  );


  buf
  g356
  (
    n441,
    n237
  );


  buf
  g357
  (
    n835,
    n309
  );


  not
  g358
  (
    n926,
    n250
  );


  not
  g359
  (
    n728,
    n290
  );


  buf
  g360
  (
    n609,
    n349
  );


  buf
  g361
  (
    n492,
    n286
  );


  not
  g362
  (
    n659,
    n221
  );


  buf
  g363
  (
    n897,
    n206
  );


  buf
  g364
  (
    n989,
    n211
  );


  not
  g365
  (
    n502,
    n194
  );


  not
  g366
  (
    n583,
    n291
  );


  not
  g367
  (
    n511,
    n323
  );


  buf
  g368
  (
    n826,
    n197
  );


  buf
  g369
  (
    n513,
    n280
  );


  buf
  g370
  (
    n551,
    n288
  );


  not
  g371
  (
    n584,
    n303
  );


  buf
  g372
  (
    n845,
    n333
  );


  buf
  g373
  (
    n660,
    n199
  );


  not
  g374
  (
    n633,
    n318
  );


  not
  g375
  (
    n642,
    n242
  );


  buf
  g376
  (
    n509,
    n277
  );


  buf
  g377
  (
    n903,
    n318
  );


  buf
  g378
  (
    n965,
    n244
  );


  not
  g379
  (
    n696,
    n292
  );


  buf
  g380
  (
    n971,
    n202
  );


  buf
  g381
  (
    n771,
    n268
  );


  buf
  g382
  (
    n671,
    n278
  );


  buf
  g383
  (
    n395,
    n213
  );


  buf
  g384
  (
    n542,
    n207
  );


  not
  g385
  (
    n425,
    n212
  );


  buf
  g386
  (
    n946,
    n340
  );


  buf
  g387
  (
    n927,
    n266
  );


  not
  g388
  (
    n378,
    n198
  );


  not
  g389
  (
    n824,
    n301
  );


  not
  g390
  (
    n808,
    n212
  );


  not
  g391
  (
    n573,
    n350
  );


  not
  g392
  (
    n442,
    n263
  );


  not
  g393
  (
    n454,
    n228
  );


  buf
  g394
  (
    n789,
    n298
  );


  buf
  g395
  (
    n383,
    n264
  );


  buf
  g396
  (
    n890,
    n289
  );


  buf
  g397
  (
    n439,
    n321
  );


  not
  g398
  (
    n577,
    n282
  );


  not
  g399
  (
    n736,
    n259
  );


  buf
  g400
  (
    n470,
    n339
  );


  buf
  g401
  (
    n924,
    n222
  );


  buf
  g402
  (
    n656,
    n243
  );


  buf
  g403
  (
    n605,
    n279
  );


  not
  g404
  (
    n475,
    n199
  );


  not
  g405
  (
    n995,
    n332
  );


  buf
  g406
  (
    n774,
    n257
  );


  not
  g407
  (
    n770,
    n243
  );


  buf
  g408
  (
    n420,
    n217
  );


  buf
  g409
  (
    n745,
    n271
  );


  buf
  g410
  (
    n777,
    n311
  );


  not
  g411
  (
    n384,
    n236
  );


  not
  g412
  (
    n374,
    n242
  );


  buf
  g413
  (
    n388,
    n260
  );


  buf
  g414
  (
    KeyWire_0_3,
    n207
  );


  not
  g415
  (
    n554,
    n338
  );


  not
  g416
  (
    n402,
    n288
  );


  not
  g417
  (
    n759,
    n240
  );


  buf
  g418
  (
    n817,
    n252
  );


  not
  g419
  (
    n920,
    n208
  );


  buf
  g420
  (
    n857,
    n269
  );


  buf
  g421
  (
    n387,
    n336
  );


  buf
  g422
  (
    n626,
    n205
  );


  not
  g423
  (
    n852,
    n274
  );


  not
  g424
  (
    n622,
    n345
  );


  buf
  g425
  (
    n486,
    n298
  );


  buf
  g426
  (
    n834,
    n234
  );


  buf
  g427
  (
    n547,
    n351
  );


  not
  g428
  (
    n459,
    n258
  );


  not
  g429
  (
    n469,
    n312
  );


  buf
  g430
  (
    n782,
    n332
  );


  buf
  g431
  (
    KeyWire_0_5,
    n200
  );


  buf
  g432
  (
    n372,
    n225
  );


  buf
  g433
  (
    n483,
    n254
  );


  buf
  g434
  (
    n401,
    n328
  );


  buf
  g435
  (
    n639,
    n281
  );


  not
  g436
  (
    n657,
    n222
  );


  buf
  g437
  (
    KeyWire_0_8,
    n326
  );


  buf
  g438
  (
    n865,
    n209
  );


  buf
  g439
  (
    n704,
    n299
  );


  buf
  g440
  (
    n977,
    n353
  );


  buf
  g441
  (
    n797,
    n319
  );


  not
  g442
  (
    n714,
    n285
  );


  not
  g443
  (
    n799,
    n346
  );


  not
  g444
  (
    n803,
    n247
  );


  buf
  g445
  (
    n467,
    n237
  );


  buf
  g446
  (
    n559,
    n282
  );


  buf
  g447
  (
    n449,
    n350
  );


  not
  g448
  (
    n781,
    n249
  );


  buf
  g449
  (
    n440,
    n259
  );


  not
  g450
  (
    n892,
    n343
  );


  buf
  g451
  (
    n679,
    n346
  );


  buf
  g452
  (
    n776,
    n232
  );


  buf
  g453
  (
    n693,
    n307
  );


  not
  g454
  (
    n804,
    n257
  );


  buf
  g455
  (
    n574,
    n230
  );


  buf
  g456
  (
    n873,
    n309
  );


  buf
  g457
  (
    n881,
    n228
  );


  not
  g458
  (
    n833,
    n241
  );


  buf
  g459
  (
    n692,
    n254
  );


  not
  g460
  (
    n686,
    n272
  );


  buf
  g461
  (
    n1001,
    n277
  );


  not
  g462
  (
    n507,
    n303
  );


  not
  g463
  (
    n739,
    n258
  );


  not
  g464
  (
    n587,
    n307
  );


  buf
  g465
  (
    n524,
    n290
  );


  buf
  g466
  (
    n592,
    n201
  );


  not
  g467
  (
    n726,
    n267
  );


  not
  g468
  (
    n641,
    n261
  );


  not
  g469
  (
    n672,
    n328
  );


  not
  g470
  (
    n687,
    n231
  );


  buf
  g471
  (
    n380,
    n218
  );


  buf
  g472
  (
    n870,
    n262
  );


  not
  g473
  (
    n405,
    n246
  );


  buf
  g474
  (
    n843,
    n214
  );


  not
  g475
  (
    n949,
    n334
  );


  not
  g476
  (
    n883,
    n224
  );


  not
  g477
  (
    n443,
    n252
  );


  not
  g478
  (
    n424,
    n335
  );


  buf
  g479
  (
    n952,
    n349
  );


  buf
  g480
  (
    n876,
    n255
  );


  not
  g481
  (
    n644,
    n221
  );


  not
  g482
  (
    n682,
    n242
  );


  not
  g483
  (
    n935,
    n261
  );


  not
  g484
  (
    n472,
    n297
  );


  not
  g485
  (
    n377,
    n317
  );


  buf
  g486
  (
    n598,
    n269
  );


  not
  g487
  (
    n539,
    n247
  );


  not
  g488
  (
    n479,
    n255
  );


  not
  g489
  (
    n512,
    n197
  );


  buf
  g490
  (
    n772,
    n327
  );


  not
  g491
  (
    n673,
    n223
  );


  not
  g492
  (
    n918,
    n229
  );


  not
  g493
  (
    n991,
    n245
  );


  buf
  g494
  (
    n900,
    n222
  );


  buf
  g495
  (
    n766,
    n288
  );


  buf
  g496
  (
    n899,
    n298
  );


  buf
  g497
  (
    n481,
    n324
  );


  buf
  g498
  (
    n861,
    n304
  );


  not
  g499
  (
    n663,
    n269
  );


  buf
  g500
  (
    n1007,
    n241
  );


  not
  g501
  (
    n731,
    n240
  );


  not
  g502
  (
    n415,
    n336
  );


  buf
  g503
  (
    n703,
    n233
  );


  buf
  g504
  (
    n600,
    n275
  );


  not
  g505
  (
    n875,
    n292
  );


  not
  g506
  (
    n879,
    n275
  );


  not
  g507
  (
    n724,
    n235
  );


  not
  g508
  (
    n521,
    n284
  );


  not
  g509
  (
    n476,
    n254
  );


  buf
  g510
  (
    n589,
    n212
  );


  buf
  g511
  (
    n794,
    n347
  );


  not
  g512
  (
    n473,
    n219
  );


  not
  g513
  (
    n893,
    n270
  );


  buf
  g514
  (
    n725,
    n322
  );


  buf
  g515
  (
    n769,
    n234
  );


  buf
  g516
  (
    n446,
    n223
  );


  buf
  g517
  (
    n910,
    n248
  );


  buf
  g518
  (
    n530,
    n202
  );


  buf
  g519
  (
    n508,
    n215
  );


  not
  g520
  (
    n968,
    n308
  );


  not
  g521
  (
    KeyWire_0_10,
    n348
  );


  buf
  g522
  (
    n668,
    n316
  );


  buf
  g523
  (
    n715,
    n265
  );


  not
  g524
  (
    n844,
    n265
  );


  not
  g525
  (
    n763,
    n332
  );


  buf
  g526
  (
    n746,
    n251
  );


  not
  g527
  (
    n718,
    n196
  );


  buf
  g528
  (
    n553,
    n227
  );


  not
  g529
  (
    n830,
    n278
  );


  buf
  g530
  (
    n477,
    n204
  );


  buf
  g531
  (
    n528,
    n295
  );


  not
  g532
  (
    n658,
    n303
  );


  not
  g533
  (
    n422,
    n330
  );


  not
  g534
  (
    n510,
    n195
  );


  buf
  g535
  (
    n563,
    n256
  );


  not
  g536
  (
    n575,
    n325
  );


  not
  g537
  (
    n818,
    n316
  );


  buf
  g538
  (
    n783,
    n308
  );


  buf
  g539
  (
    n964,
    n338
  );


  not
  g540
  (
    n677,
    n330
  );


  buf
  g541
  (
    n1008,
    n310
  );


  buf
  g542
  (
    n755,
    n329
  );


  buf
  g543
  (
    n576,
    n295
  );


  not
  g544
  (
    n571,
    n345
  );


  buf
  g545
  (
    n406,
    n292
  );


  not
  g546
  (
    n485,
    n270
  );


  buf
  g547
  (
    n458,
    n247
  );


  not
  g548
  (
    n992,
    n282
  );


  buf
  g549
  (
    n859,
    n271
  );


  buf
  g550
  (
    n988,
    n343
  );


  buf
  g551
  (
    n921,
    n352
  );


  not
  g552
  (
    n842,
    n196
  );


  buf
  g553
  (
    n675,
    n248
  );


  buf
  g554
  (
    n711,
    n281
  );


  buf
  g555
  (
    n868,
    n212
  );


  buf
  g556
  (
    n912,
    n274
  );


  not
  g557
  (
    n465,
    n352
  );


  buf
  g558
  (
    n1000,
    n339
  );


  buf
  g559
  (
    n582,
    n283
  );


  buf
  g560
  (
    n670,
    n225
  );


  not
  g561
  (
    n588,
    n238
  );


  not
  g562
  (
    n594,
    n309
  );


  buf
  g563
  (
    n389,
    n314
  );


  not
  g564
  (
    n408,
    n268
  );


  buf
  g565
  (
    n878,
    n325
  );


  not
  g566
  (
    n778,
    n323
  );


  not
  g567
  (
    n815,
    n337
  );


  not
  g568
  (
    n945,
    n353
  );


  buf
  g569
  (
    n555,
    n235
  );


  buf
  g570
  (
    n557,
    n263
  );


  not
  g571
  (
    n394,
    n296
  );


  not
  g572
  (
    n690,
    n279
  );


  buf
  g573
  (
    n515,
    n277
  );


  buf
  g574
  (
    n496,
    n280
  );


  not
  g575
  (
    n618,
    n331
  );


  not
  g576
  (
    n386,
    n233
  );


  buf
  g577
  (
    n955,
    n350
  );


  buf
  g578
  (
    n923,
    n351
  );


  not
  g579
  (
    n450,
    n344
  );


  buf
  g580
  (
    n471,
    n210
  );


  buf
  g581
  (
    n966,
    n221
  );


  not
  g582
  (
    n651,
    n216
  );


  buf
  g583
  (
    n733,
    n294
  );


  buf
  g584
  (
    n747,
    n211
  );


  not
  g585
  (
    n649,
    n253
  );


  not
  g586
  (
    n620,
    n200
  );


  buf
  g587
  (
    n560,
    n215
  );


  buf
  g588
  (
    n706,
    n198
  );


  buf
  g589
  (
    n438,
    n244
  );


  not
  g590
  (
    n712,
    n233
  );


  buf
  g591
  (
    n790,
    n220
  );


  buf
  g592
  (
    n648,
    n335
  );


  not
  g593
  (
    n957,
    n309
  );


  buf
  g594
  (
    n810,
    n240
  );


  buf
  g595
  (
    n956,
    n267
  );


  buf
  g596
  (
    n943,
    n260
  );


  buf
  g597
  (
    n652,
    n224
  );


  not
  g598
  (
    n902,
    n238
  );


  not
  g599
  (
    n788,
    n226
  );


  buf
  g600
  (
    n540,
    n301
  );


  not
  g601
  (
    n872,
    n231
  );


  not
  g602
  (
    n831,
    n310
  );


  not
  g603
  (
    n742,
    n297
  );


  not
  g604
  (
    n697,
    n275
  );


  buf
  g605
  (
    n727,
    n285
  );


  not
  g606
  (
    n904,
    n331
  );


  not
  g607
  (
    n860,
    n349
  );


  not
  g608
  (
    n457,
    n257
  );


  not
  g609
  (
    n534,
    n342
  );


  buf
  g610
  (
    n767,
    n196
  );


  buf
  g611
  (
    n619,
    n206
  );


  not
  g612
  (
    n432,
    n200
  );


  not
  g613
  (
    n517,
    n332
  );


  not
  g614
  (
    KeyWire_0_0,
    n299
  );


  buf
  g615
  (
    n461,
    n338
  );


  buf
  g616
  (
    n825,
    n249
  );


  not
  g617
  (
    n417,
    n229
  );


  not
  g618
  (
    n722,
    n242
  );


  buf
  g619
  (
    n667,
    n263
  );


  not
  g620
  (
    n578,
    n248
  );


  buf
  g621
  (
    n421,
    n230
  );


  buf
  g622
  (
    n418,
    n302
  );


  buf
  g623
  (
    n669,
    n232
  );


  buf
  g624
  (
    n579,
    n194
  );


  buf
  g625
  (
    n445,
    n207
  );


  buf
  g626
  (
    n428,
    n271
  );


  buf
  g627
  (
    n640,
    n341
  );


  buf
  g628
  (
    n664,
    n252
  );


  not
  g629
  (
    n779,
    n305
  );


  not
  g630
  (
    n716,
    n236
  );


  buf
  g631
  (
    n986,
    n246
  );


  buf
  g632
  (
    n828,
    n294
  );


  not
  g633
  (
    n552,
    n278
  );


  not
  g634
  (
    n916,
    n220
  );


  not
  g635
  (
    n849,
    n342
  );


  buf
  g636
  (
    n764,
    n217
  );


  not
  g637
  (
    n630,
    n265
  );


  buf
  g638
  (
    n546,
    n256
  );


  not
  g639
  (
    n397,
    n295
  );


  not
  g640
  (
    n780,
    n281
  );


  not
  g641
  (
    n953,
    n310
  );


  buf
  g642
  (
    n967,
    n223
  );


  not
  g643
  (
    n795,
    n334
  );


  not
  g644
  (
    n846,
    n223
  );


  not
  g645
  (
    n898,
    n283
  );


  buf
  g646
  (
    n911,
    n315
  );


  not
  g647
  (
    n678,
    n220
  );


  not
  g648
  (
    n720,
    n290
  );


  buf
  g649
  (
    n909,
    n310
  );


  buf
  g650
  (
    n942,
    n322
  );


  buf
  g651
  (
    n694,
    n220
  );


  not
  g652
  (
    n604,
    n213
  );


  not
  g653
  (
    n832,
    n329
  );


  buf
  g654
  (
    n951,
    n335
  );


  not
  g655
  (
    n922,
    n320
  );


  not
  g656
  (
    n721,
    n218
  );


  buf
  g657
  (
    n959,
    n337
  );


  not
  g658
  (
    n984,
    n219
  );


  buf
  g659
  (
    n556,
    n245
  );


  not
  g660
  (
    n816,
    n304
  );


  buf
  g661
  (
    n568,
    n248
  );


  buf
  g662
  (
    KeyWire_0_1,
    n300
  );


  buf
  g663
  (
    n997,
    n251
  );


  not
  g664
  (
    n885,
    n284
  );


  not
  g665
  (
    n787,
    n313
  );


  not
  g666
  (
    n925,
    n273
  );


  buf
  g667
  (
    n896,
    n287
  );


  not
  g668
  (
    n735,
    n246
  );


  not
  g669
  (
    n891,
    n199
  );


  buf
  g670
  (
    n504,
    n258
  );


  buf
  g671
  (
    n653,
    n256
  );


  buf
  g672
  (
    n529,
    n255
  );


  not
  g673
  (
    n681,
    n320
  );


  not
  g674
  (
    n647,
    n350
  );


  not
  g675
  (
    n646,
    n340
  );


  not
  g676
  (
    n806,
    n285
  );


  buf
  g677
  (
    n732,
    n308
  );


  not
  g678
  (
    n848,
    n308
  );


  not
  g679
  (
    n749,
    n298
  );


  not
  g680
  (
    n490,
    n311
  );


  not
  g681
  (
    n596,
    n194
  );


  buf
  g682
  (
    n550,
    n227
  );


  not
  g683
  (
    n456,
    n246
  );


  not
  g684
  (
    n569,
    n317
  );


  not
  g685
  (
    n423,
    n206
  );


  buf
  g686
  (
    n506,
    n326
  );


  buf
  g687
  (
    n635,
    n293
  );


  buf
  g688
  (
    n612,
    n304
  );


  buf
  g689
  (
    n409,
    n333
  );


  buf
  g690
  (
    n753,
    n241
  );


  buf
  g691
  (
    n887,
    n262
  );


  not
  g692
  (
    n981,
    n268
  );


  not
  g693
  (
    n522,
    n239
  );


  not
  g694
  (
    n978,
    n289
  );


  buf
  g695
  (
    n938,
    n261
  );


  buf
  g696
  (
    n708,
    n209
  );


  not
  g697
  (
    n480,
    n270
  );


  not
  g698
  (
    n468,
    n342
  );


  not
  g699
  (
    n980,
    n268
  );


  not
  g700
  (
    n814,
    n293
  );


  buf
  g701
  (
    n602,
    n333
  );


  not
  g702
  (
    n549,
    n203
  );


  not
  g703
  (
    n381,
    n351
  );


  buf
  g704
  (
    n614,
    n211
  );


  not
  g705
  (
    n932,
    n283
  );


  buf
  g706
  (
    n734,
    n235
  );


  buf
  g707
  (
    n391,
    n213
  );


  not
  g708
  (
    n717,
    n222
  );


  buf
  g709
  (
    n562,
    n228
  );


  not
  g710
  (
    n974,
    n210
  );


  buf
  g711
  (
    n838,
    n226
  );


  not
  g712
  (
    n497,
    n211
  );


  buf
  g713
  (
    n983,
    n265
  );


  not
  g714
  (
    n785,
    n291
  );


  not
  g715
  (
    n413,
    n208
  );


  not
  g716
  (
    n866,
    n214
  );


  buf
  g717
  (
    n464,
    n337
  );


  buf
  g718
  (
    n548,
    n322
  );


  not
  g719
  (
    n453,
    n259
  );


  not
  g720
  (
    n869,
    n336
  );


  buf
  g721
  (
    n793,
    n280
  );


  buf
  g722
  (
    n393,
    n299
  );


  not
  g723
  (
    n707,
    n255
  );


  not
  g724
  (
    n437,
    n329
  );


  not
  g725
  (
    KeyWire_0_11,
    n195
  );


  not
  g726
  (
    n863,
    n273
  );


  not
  g727
  (
    n796,
    n347
  );


  buf
  g728
  (
    n392,
    n315
  );


  buf
  g729
  (
    n856,
    n197
  );


  buf
  g730
  (
    n705,
    n307
  );


  buf
  g731
  (
    n930,
    n226
  );


  buf
  g732
  (
    n894,
    n297
  );


  not
  g733
  (
    n954,
    n272
  );


  not
  g734
  (
    n533,
    n284
  );


  buf
  g735
  (
    n370,
    n325
  );


  buf
  g736
  (
    n855,
    n327
  );


  not
  g737
  (
    n979,
    n296
  );


  not
  g738
  (
    n403,
    n289
  );


  buf
  g739
  (
    n400,
    n235
  );


  buf
  g740
  (
    n572,
    n318
  );


  buf
  g741
  (
    n928,
    n216
  );


  not
  g742
  (
    n654,
    n225
  );


  not
  g743
  (
    n590,
    n203
  );


  not
  g744
  (
    n434,
    n218
  );


  not
  g745
  (
    n754,
    n348
  );


  buf
  g746
  (
    n915,
    n239
  );


  not
  g747
  (
    n623,
    n286
  );


  buf
  g748
  (
    n791,
    n294
  );


  buf
  g749
  (
    n829,
    n352
  );


  buf
  g750
  (
    n827,
    n205
  );


  buf
  g751
  (
    n994,
    n272
  );


  not
  g752
  (
    n934,
    n210
  );


  not
  g753
  (
    n518,
    n294
  );


  not
  g754
  (
    n895,
    n324
  );


  buf
  g755
  (
    n792,
    n245
  );


  buf
  g756
  (
    n773,
    n249
  );


  buf
  g757
  (
    n411,
    n351
  );


  not
  g758
  (
    n751,
    n343
  );


  not
  g759
  (
    n611,
    n291
  );


  not
  g760
  (
    n455,
    n339
  );


  buf
  g761
  (
    n823,
    n300
  );


  buf
  g762
  (
    n631,
    n195
  );


  buf
  g763
  (
    n836,
    n278
  );


  buf
  g764
  (
    n689,
    n206
  );


  buf
  g765
  (
    n740,
    n326
  );


  not
  g766
  (
    n847,
    n347
  );


  buf
  g767
  (
    n608,
    n295
  );


  not
  g768
  (
    n1006,
    n347
  );


  not
  g769
  (
    n990,
    n208
  );


  not
  g770
  (
    n801,
    n346
  );


  buf
  g771
  (
    n937,
    n341
  );


  buf
  g772
  (
    n882,
    n203
  );


  buf
  g773
  (
    n595,
    n236
  );


  not
  g774
  (
    n864,
    n276
  );


  not
  g775
  (
    n744,
    n244
  );


  not
  g776
  (
    n812,
    n213
  );


  not
  g777
  (
    n889,
    n341
  );


  not
  g778
  (
    n474,
    n217
  );


  buf
  g779
  (
    n858,
    n305
  );


  buf
  g780
  (
    n613,
    n219
  );


  buf
  g781
  (
    n680,
    n313
  );


  not
  g782
  (
    n503,
    n197
  );


  buf
  g783
  (
    n385,
    n287
  );


  not
  g784
  (
    n960,
    n209
  );


  buf
  g785
  (
    n514,
    n293
  );


  not
  g786
  (
    n581,
    n302
  );


  buf
  g787
  (
    n699,
    n238
  );


  not
  g788
  (
    n650,
    n217
  );


  buf
  g789
  (
    n975,
    n288
  );


  not
  g790
  (
    KeyWire_0_7,
    n313
  );


  buf
  g791
  (
    n813,
    n352
  );


  not
  g792
  (
    n839,
    n216
  );


  buf
  g793
  (
    n743,
    n317
  );


  not
  g794
  (
    n632,
    n279
  );


  not
  g795
  (
    n625,
    n273
  );


  buf
  g796
  (
    n629,
    n199
  );


  buf
  g797
  (
    n536,
    n215
  );


  buf
  g798
  (
    n525,
    n272
  );


  buf
  g799
  (
    KeyWire_0_6,
    n344
  );


  buf
  g800
  (
    n390,
    n348
  );


  buf
  g801
  (
    n585,
    n296
  );


  buf
  g802
  (
    n463,
    n250
  );


  buf
  g803
  (
    n800,
    n262
  );


  not
  g804
  (
    n607,
    n236
  );


  buf
  g805
  (
    n558,
    n346
  );


  not
  g806
  (
    n939,
    n252
  );


  not
  g807
  (
    n535,
    n321
  );


  buf
  g808
  (
    n821,
    n202
  );


  not
  g809
  (
    n752,
    n345
  );


  buf
  g810
  (
    n435,
    n311
  );


  buf
  g811
  (
    n987,
    n227
  );


  buf
  g812
  (
    n691,
    n323
  );


  not
  g813
  (
    n580,
    n237
  );


  buf
  g814
  (
    n488,
    n301
  );


  not
  g815
  (
    n599,
    n344
  );


  not
  g816
  (
    n805,
    n286
  );


  not
  g817
  (
    n570,
    n266
  );


  not
  g818
  (
    n917,
    n230
  );


  not
  g819
  (
    n985,
    n340
  );


  buf
  g820
  (
    n685,
    n296
  );


  buf
  g821
  (
    n820,
    n329
  );


  buf
  g822
  (
    n505,
    n343
  );


  buf
  g823
  (
    n634,
    n202
  );


  not
  g824
  (
    n907,
    n312
  );


  not
  g825
  (
    n982,
    n312
  );


  buf
  g826
  (
    n841,
    n324
  );


  not
  g827
  (
    n615,
    n239
  );


  not
  g828
  (
    n527,
    n335
  );


  not
  g829
  (
    n436,
    n214
  );


  buf
  g830
  (
    n482,
    n306
  );


  buf
  g831
  (
    n655,
    n259
  );


  not
  g832
  (
    n962,
    n210
  );


  not
  g833
  (
    n947,
    n302
  );


  buf
  g834
  (
    n809,
    n276
  );


  not
  g835
  (
    n447,
    n232
  );


  buf
  g836
  (
    n802,
    n330
  );


  not
  g837
  (
    n407,
    n304
  );


  not
  g838
  (
    n944,
    n312
  );


  not
  g839
  (
    n948,
    n205
  );


  buf
  g840
  (
    n741,
    n253
  );


  buf
  g841
  (
    n901,
    n232
  );


  buf
  g842
  (
    n462,
    n336
  );


  not
  g843
  (
    n698,
    n234
  );


  buf
  g844
  (
    n666,
    n275
  );


  not
  g845
  (
    n494,
    n225
  );


  buf
  g846
  (
    n586,
    n306
  );


  buf
  g847
  (
    n760,
    n201
  );


  not
  g848
  (
    n451,
    n293
  );


  not
  g849
  (
    n601,
    n306
  );


  buf
  g850
  (
    n498,
    n234
  );


  buf
  g851
  (
    n963,
    n319
  );


  not
  g852
  (
    n906,
    n301
  );


  not
  g853
  (
    n913,
    n284
  );


  not
  g854
  (
    n1004,
    n340
  );


  buf
  g855
  (
    n683,
    n271
  );


  not
  g856
  (
    n404,
    n315
  );


  buf
  g857
  (
    n702,
    n264
  );


  buf
  g858
  (
    n516,
    n203
  );


  not
  g859
  (
    n684,
    n243
  );


  not
  g860
  (
    n936,
    n269
  );


  buf
  g861
  (
    n853,
    n324
  );


  not
  g862
  (
    n501,
    n226
  );


  buf
  g863
  (
    n940,
    n313
  );


  buf
  g864
  (
    n564,
    n237
  );


  not
  g865
  (
    n567,
    n321
  );


  buf
  g866
  (
    n561,
    n349
  );


  buf
  g867
  (
    n757,
    n266
  );


  buf
  g868
  (
    n961,
    n334
  );


  buf
  g869
  (
    n996,
    n198
  );


  buf
  g870
  (
    n532,
    n307
  );


  buf
  g871
  (
    n636,
    n302
  );


  buf
  g872
  (
    n886,
    n227
  );


  not
  g873
  (
    n478,
    n353
  );


  not
  g874
  (
    n376,
    n256
  );


  not
  g875
  (
    n854,
    n327
  );


  buf
  g876
  (
    n972,
    n264
  );


  not
  g877
  (
    n695,
    n291
  );


  not
  g878
  (
    n908,
    n345
  );


  buf
  g879
  (
    n637,
    n274
  );


  not
  g880
  (
    n621,
    n322
  );


  buf
  g881
  (
    n427,
    n270
  );


  buf
  g882
  (
    n768,
    n321
  );


  buf
  g883
  (
    n610,
    n238
  );


  not
  g884
  (
    n375,
    n253
  );


  not
  g885
  (
    n628,
    n344
  );


  not
  g886
  (
    n998,
    n315
  );


  not
  g887
  (
    n373,
    n208
  );


  buf
  g888
  (
    n862,
    n201
  );


  buf
  g889
  (
    n627,
    n300
  );


  buf
  g890
  (
    n969,
    n276
  );


  not
  g891
  (
    n448,
    n286
  );


  not
  g892
  (
    n941,
    n300
  );


  not
  g893
  (
    n676,
    n224
  );


  buf
  g894
  (
    n877,
    n326
  );


  buf
  g895
  (
    n412,
    n251
  );


  not
  g896
  (
    n765,
    n334
  );


  not
  g897
  (
    n784,
    n281
  );


  not
  g898
  (
    n500,
    n306
  );


  buf
  g899
  (
    n688,
    n253
  );


  buf
  g900
  (
    n460,
    n325
  );


  buf
  g901
  (
    n371,
    n285
  );


  not
  g902
  (
    n444,
    n330
  );


  not
  g903
  (
    n958,
    n314
  );


  not
  g904
  (
    n874,
    n229
  );


  not
  g905
  (
    n487,
    n318
  );


  buf
  g906
  (
    n761,
    n221
  );


  buf
  g907
  (
    n526,
    n204
  );


  not
  g908
  (
    n674,
    n230
  );


  buf
  g909
  (
    n543,
    n266
  );


  not
  g910
  (
    n491,
    n314
  );


  buf
  g911
  (
    n884,
    n204
  );


  buf
  g912
  (
    n710,
    n201
  );


  not
  g913
  (
    n850,
    n207
  );


  not
  g914
  (
    n643,
    n247
  );


  buf
  g915
  (
    n871,
    n264
  );


  not
  g916
  (
    n933,
    n267
  );


  buf
  g917
  (
    n737,
    n233
  );


  not
  g918
  (
    n762,
    n338
  );


  buf
  g919
  (
    n538,
    n244
  );


  buf
  g920
  (
    n606,
    n323
  );


  not
  g921
  (
    n786,
    n280
  );


  buf
  g922
  (
    n545,
    n245
  );


  not
  g923
  (
    n419,
    n274
  );


  not
  g924
  (
    n700,
    n204
  );


  not
  g925
  (
    n709,
    n215
  );


  buf
  g926
  (
    n489,
    n311
  );


  not
  g927
  (
    n398,
    n195
  );


  not
  g928
  (
    n819,
    n254
  );


  buf
  g929
  (
    n851,
    n194
  );


  buf
  g930
  (
    n399,
    n290
  );


  not
  g931
  (
    n807,
    n277
  );


  buf
  g932
  (
    n379,
    n283
  );


  buf
  g933
  (
    n905,
    n328
  );


  buf
  g934
  (
    n414,
    n249
  );


  buf
  g935
  (
    n811,
    n314
  );


  buf
  g936
  (
    n822,
    n216
  );


  buf
  g937
  (
    n661,
    n258
  );


  buf
  g938
  (
    n758,
    n263
  );


  buf
  g939
  (
    n433,
    n331
  );


  not
  g940
  (
    n499,
    n243
  );


  buf
  g941
  (
    n662,
    n282
  );


  buf
  g942
  (
    n888,
    n228
  );


  not
  g943
  (
    n730,
    n348
  );


  not
  g944
  (
    n616,
    n316
  );


  buf
  g945
  (
    n976,
    n305
  );


  buf
  g946
  (
    n929,
    n305
  );


  not
  g947
  (
    n531,
    n240
  );


  not
  g948
  (
    n665,
    n262
  );


  not
  g949
  (
    n519,
    n260
  );


  buf
  g950
  (
    n645,
    n331
  );


  not
  g951
  (
    n867,
    n297
  );


  not
  g952
  (
    n719,
    n219
  );


  buf
  g953
  (
    n931,
    n239
  );


  buf
  g954
  (
    n1003,
    n209
  );


  not
  g955
  (
    n410,
    n316
  );


  buf
  g956
  (
    n565,
    n279
  );


  not
  g957
  (
    n382,
    n231
  );


  not
  g958
  (
    n1002,
    n289
  );


  not
  g959
  (
    n431,
    n218
  );


  buf
  g960
  (
    n919,
    n276
  );


  not
  g961
  (
    n914,
    n224
  );


  buf
  g962
  (
    n999,
    n320
  );


  not
  g963
  (
    n523,
    n250
  );


  not
  g964
  (
    n756,
    n320
  );


  not
  g965
  (
    n429,
    n251
  );


  not
  g966
  (
    n396,
    n260
  );


  not
  g967
  (
    n701,
    n261
  );


  buf
  g968
  (
    n738,
    n287
  );


  not
  g969
  (
    n970,
    n241
  );


  not
  g970
  (
    n775,
    n229
  );


  not
  g971
  (
    n597,
    n341
  );


  buf
  g972
  (
    n495,
    n299
  );


  buf
  g973
  (
    n729,
    n303
  );


  buf
  g974
  (
    n603,
    n231
  );


  not
  g975
  (
    n537,
    n273
  );


  nor
  g976
  (
    n1484,
    n674,
    n392,
    n774,
    n890
  );


  xnor
  g977
  (
    n1210,
    n584,
    n917,
    n669,
    n608
  );


  nand
  g978
  (
    n1032,
    n511,
    n733,
    n612,
    n843
  );


  nor
  g979
  (
    n1209,
    n897,
    n870,
    n539,
    n730
  );


  xnor
  g980
  (
    n1274,
    n956,
    n773,
    n681,
    n490
  );


  and
  g981
  (
    n1559,
    n973,
    n448,
    n751,
    n596
  );


  and
  g982
  (
    n1169,
    n783,
    n521,
    n893,
    n814
  );


  nor
  g983
  (
    n1340,
    n845,
    n551,
    n514,
    n438
  );


  nor
  g984
  (
    n1354,
    n582,
    n703,
    n739,
    n777
  );


  and
  g985
  (
    n1299,
    n491,
    n803,
    n967,
    n562
  );


  xor
  g986
  (
    n1279,
    n418,
    n688,
    n837,
    n700
  );


  or
  g987
  (
    n1157,
    n453,
    n606,
    n971,
    n545
  );


  nor
  g988
  (
    n1261,
    n606,
    n929,
    n820,
    n790
  );


  xnor
  g989
  (
    n1113,
    n601,
    n739,
    n790,
    n799
  );


  and
  g990
  (
    n1557,
    n661,
    n729,
    n711,
    n859
  );


  or
  g991
  (
    n1234,
    n899,
    n784,
    n574,
    n680
  );


  xnor
  g992
  (
    n1516,
    n811,
    n500,
    n875,
    n542
  );


  xnor
  g993
  (
    n1416,
    n778,
    n941,
    n656,
    n494
  );


  xor
  g994
  (
    n1486,
    n485,
    n482,
    n798,
    n816
  );


  xnor
  g995
  (
    n1370,
    n621,
    n742,
    n877,
    n909
  );


  xor
  g996
  (
    n1170,
    n849,
    n446,
    n608,
    n837
  );


  xor
  g997
  (
    n1499,
    n602,
    n592,
    n572,
    n588
  );


  nand
  g998
  (
    n1237,
    n892,
    n560,
    n885,
    n715
  );


  nor
  g999
  (
    n1342,
    n516,
    n782,
    n402,
    n818
  );


  and
  g1000
  (
    n1387,
    n983,
    n698,
    n965,
    n744
  );


  xnor
  g1001
  (
    n1211,
    n552,
    n378,
    n903,
    n676
  );


  nand
  g1002
  (
    n1217,
    n685,
    n896,
    n484,
    n629
  );


  or
  g1003
  (
    n1052,
    n507,
    n823,
    n672,
    n695
  );


  nand
  g1004
  (
    n1351,
    n623,
    n634,
    n596,
    n938
  );


  nand
  g1005
  (
    n1242,
    n528,
    n519,
    n716,
    n523
  );


  and
  g1006
  (
    n1336,
    n471,
    n871,
    n832,
    n597
  );


  xor
  g1007
  (
    n1412,
    n656,
    n841,
    n509,
    n519
  );


  xnor
  g1008
  (
    n1284,
    n819,
    n470,
    n810,
    n866
  );


  nor
  g1009
  (
    n1315,
    n443,
    n934,
    n807,
    n604
  );


  nor
  g1010
  (
    n1158,
    n862,
    n973,
    n639,
    n859
  );


  xnor
  g1011
  (
    n1436,
    n537,
    n812,
    n822,
    n986
  );


  xor
  g1012
  (
    n1467,
    n809,
    n793,
    n840,
    n973
  );


  nand
  g1013
  (
    n1479,
    n858,
    n680,
    n779,
    n386
  );


  xor
  g1014
  (
    n1422,
    n805,
    n886,
    n392,
    n954
  );


  nor
  g1015
  (
    n1087,
    n686,
    n828,
    n722,
    n454
  );


  and
  g1016
  (
    n1365,
    n458,
    n953,
    n973,
    n664
  );


  xor
  g1017
  (
    n1045,
    n476,
    n476,
    n537,
    n829
  );


  or
  g1018
  (
    n1439,
    n426,
    n988,
    n961,
    n842
  );


  nor
  g1019
  (
    n1154,
    n912,
    n932,
    n727,
    n663
  );


  nor
  g1020
  (
    n1190,
    n507,
    n745,
    n545,
    n461
  );


  xnor
  g1021
  (
    n1017,
    n618,
    n717,
    n817,
    n828
  );


  and
  g1022
  (
    n1377,
    n735,
    n612,
    n434,
    n817
  );


  or
  g1023
  (
    n1084,
    n955,
    n945,
    n585,
    n494
  );


  xnor
  g1024
  (
    n1325,
    n789,
    n468,
    n844,
    n882
  );


  nor
  g1025
  (
    n1569,
    n936,
    n748,
    n483,
    n591
  );


  and
  g1026
  (
    n1163,
    n722,
    n783,
    n532,
    n643
  );


  xnor
  g1027
  (
    n1303,
    n985,
    n897,
    n861,
    n755
  );


  nand
  g1028
  (
    n1395,
    n796,
    n980,
    n810,
    n409
  );


  xor
  g1029
  (
    n1366,
    n393,
    n464,
    n714,
    n825
  );


  or
  g1030
  (
    n1291,
    n758,
    n792,
    n633,
    n910
  );


  and
  g1031
  (
    n1264,
    n800,
    n551,
    n646,
    n979
  );


  nand
  g1032
  (
    n1272,
    n679,
    n571,
    n594,
    n766
  );


  and
  g1033
  (
    n1310,
    n920,
    n730,
    n855,
    n970
  );


  nor
  g1034
  (
    n1500,
    n981,
    n516,
    n966,
    n387
  );


  or
  g1035
  (
    n1584,
    n909,
    n655,
    n857,
    n615
  );


  and
  g1036
  (
    n1253,
    n467,
    n461,
    n546,
    n864
  );


  or
  g1037
  (
    n1587,
    n610,
    n419,
    n773,
    n467
  );


  nor
  g1038
  (
    n1060,
    n788,
    n515,
    n716,
    n746
  );


  nand
  g1039
  (
    n1225,
    n661,
    n982,
    n863,
    n964
  );


  or
  g1040
  (
    n1320,
    n696,
    n938,
    n776,
    n385
  );


  nor
  g1041
  (
    n1596,
    n550,
    n814,
    n900,
    n876
  );


  xor
  g1042
  (
    n1555,
    n704,
    n605,
    n661,
    n719
  );


  xor
  g1043
  (
    n1338,
    n713,
    n702,
    n671,
    n657
  );


  nor
  g1044
  (
    n1227,
    n416,
    n480,
    n905,
    n486
  );


  and
  g1045
  (
    n1179,
    n534,
    n914,
    n920,
    n946
  );


  xnor
  g1046
  (
    n1203,
    n632,
    n830,
    n503,
    n979
  );


  or
  g1047
  (
    n1355,
    n611,
    n551,
    n830,
    n554
  );


  nor
  g1048
  (
    n1498,
    n906,
    n561,
    n741,
    n539
  );


  xnor
  g1049
  (
    n1330,
    n579,
    n823,
    n802,
    n615
  );


  xnor
  g1050
  (
    n1260,
    n849,
    n481,
    n895,
    n718
  );


  nand
  g1051
  (
    n1438,
    n492,
    n569,
    n980,
    n682
  );


  xnor
  g1052
  (
    n1404,
    n734,
    n486,
    n617,
    n753
  );


  and
  g1053
  (
    n1509,
    n943,
    n950,
    n878,
    n645
  );


  and
  g1054
  (
    n1530,
    n437,
    n750,
    n732,
    n411
  );


  xor
  g1055
  (
    n1181,
    n567,
    n451,
    n487,
    n775
  );


  or
  g1056
  (
    n1413,
    n822,
    n587,
    n813,
    n869
  );


  xor
  g1057
  (
    n1139,
    n469,
    n789,
    n600,
    n728
  );


  and
  g1058
  (
    n1111,
    n471,
    n549,
    n750,
    n660
  );


  xor
  g1059
  (
    n1164,
    n754,
    n626,
    n923,
    n526
  );


  xnor
  g1060
  (
    n1257,
    n592,
    n490,
    n586,
    n860
  );


  and
  g1061
  (
    n1301,
    n932,
    n537,
    n479,
    n706
  );


  nor
  g1062
  (
    n1361,
    n732,
    n564,
    n529,
    n476
  );


  or
  g1063
  (
    n1363,
    n950,
    n681,
    n541,
    n888
  );


  xor
  g1064
  (
    n1477,
    n657,
    n556,
    n862,
    n752
  );


  or
  g1065
  (
    n1451,
    n770,
    n790,
    n699,
    n712
  );


  xor
  g1066
  (
    n1490,
    n571,
    n667,
    n457,
    n597
  );


  xor
  g1067
  (
    n1251,
    n899,
    n509,
    n958,
    n598
  );


  xor
  g1068
  (
    n1463,
    n880,
    n473,
    n812,
    n956
  );


  or
  g1069
  (
    n1398,
    n922,
    n959,
    n450,
    n936
  );


  xor
  g1070
  (
    n1040,
    n879,
    n987,
    n945,
    n685
  );


  and
  g1071
  (
    n1376,
    n845,
    n492,
    n744,
    n710
  );


  and
  g1072
  (
    n1537,
    n603,
    n659,
    n700,
    n746
  );


  nand
  g1073
  (
    n1380,
    n785,
    n770,
    n462,
    n848
  );


  nand
  g1074
  (
    n1345,
    n620,
    n564,
    n413,
    n417
  );


  or
  g1075
  (
    n1042,
    n943,
    n894,
    n799,
    n837
  );


  and
  g1076
  (
    n1071,
    n622,
    n939,
    n540,
    n797
  );


  and
  g1077
  (
    n1184,
    n879,
    n749,
    n502,
    n519
  );


  or
  g1078
  (
    n1137,
    n864,
    n517,
    n429,
    n989
  );


  xnor
  g1079
  (
    n1200,
    n422,
    n933,
    n431,
    n860
  );


  or
  g1080
  (
    n1009,
    n573,
    n477,
    n534,
    n374
  );


  nand
  g1081
  (
    n1570,
    n535,
    n959,
    n968,
    n636
  );


  and
  g1082
  (
    n1494,
    n709,
    n878,
    n487,
    n977
  );


  nor
  g1083
  (
    n1344,
    n522,
    n595,
    n795,
    n821
  );


  xnor
  g1084
  (
    n1464,
    n964,
    n454,
    n425,
    n717
  );


  or
  g1085
  (
    n1278,
    n599,
    n649,
    n661,
    n916
  );


  and
  g1086
  (
    n1214,
    n428,
    n620,
    n715,
    n498
  );


  and
  g1087
  (
    n1597,
    n621,
    n394,
    n967,
    n719
  );


  or
  g1088
  (
    n1024,
    n582,
    n737,
    n465,
    n850
  );


  nor
  g1089
  (
    n1396,
    n414,
    n614,
    n427,
    n940
  );


  or
  g1090
  (
    n1048,
    n574,
    n639,
    n627,
    n426
  );


  nor
  g1091
  (
    n1240,
    n527,
    n563,
    n491,
    n532
  );


  or
  g1092
  (
    n1583,
    n597,
    n533,
    n735,
    n499
  );


  or
  g1093
  (
    n1580,
    n435,
    n931,
    n442,
    n437
  );


  nor
  g1094
  (
    n1304,
    n806,
    n379,
    n626,
    n452
  );


  or
  g1095
  (
    n1527,
    n862,
    n444,
    n642,
    n740
  );


  or
  g1096
  (
    n1456,
    n726,
    n642,
    n754,
    n915
  );


  nor
  g1097
  (
    n1465,
    n450,
    n602,
    n667,
    n726
  );


  or
  g1098
  (
    n1382,
    n410,
    n835,
    n557,
    n521
  );


  and
  g1099
  (
    n1318,
    n787,
    n986,
    n511,
    n453
  );


  xor
  g1100
  (
    n1302,
    n752,
    n688,
    n765,
    n666
  );


  xnor
  g1101
  (
    n1452,
    n719,
    n460,
    n813,
    n703
  );


  xor
  g1102
  (
    n1187,
    n442,
    n613,
    n731,
    n670
  );


  xor
  g1103
  (
    n1512,
    n690,
    n772,
    n851,
    n491
  );


  and
  g1104
  (
    n1089,
    n689,
    n613,
    n656,
    n424
  );


  nor
  g1105
  (
    n1534,
    n797,
    n547,
    n485,
    n789
  );


  xor
  g1106
  (
    n1255,
    n579,
    n609,
    n455,
    n720
  );


  nor
  g1107
  (
    n1079,
    n972,
    n652,
    n739,
    n662
  );


  nand
  g1108
  (
    n1492,
    n639,
    n675,
    n577,
    n801
  );


  and
  g1109
  (
    KeyWire_0_12,
    n963,
    n794,
    n917,
    n476
  );


  nand
  g1110
  (
    n1189,
    n609,
    n569,
    n958,
    n819
  );


  nand
  g1111
  (
    n1077,
    n727,
    n658,
    n677,
    n607
  );


  xor
  g1112
  (
    n1081,
    n385,
    n554,
    n750,
    n429
  );


  nor
  g1113
  (
    n1522,
    n882,
    n894,
    n933,
    n598
  );


  and
  g1114
  (
    n1589,
    n560,
    n795,
    n683,
    n747
  );


  xnor
  g1115
  (
    n1473,
    n782,
    n692,
    n478,
    n496
  );


  nor
  g1116
  (
    n1120,
    n870,
    n664,
    n463,
    n758
  );


  and
  g1117
  (
    n1035,
    n859,
    n905,
    n536,
    n625
  );


  or
  g1118
  (
    n1581,
    n445,
    n721,
    n425,
    n552
  );


  nand
  g1119
  (
    n1127,
    n512,
    n581,
    n398,
    n723
  );


  xor
  g1120
  (
    n1266,
    n497,
    n975,
    n905,
    n600
  );


  xor
  g1121
  (
    n1461,
    n946,
    n904,
    n873,
    n456
  );


  nand
  g1122
  (
    n1028,
    n585,
    n714,
    n724,
    n902
  );


  xnor
  g1123
  (
    n1540,
    n594,
    n624,
    n578,
    n711
  );


  nand
  g1124
  (
    n1076,
    n831,
    n878,
    n593,
    n570
  );


  nand
  g1125
  (
    n1142,
    n887,
    n559,
    n964,
    n716
  );


  nor
  g1126
  (
    n1223,
    n493,
    n512,
    n578,
    n695
  );


  or
  g1127
  (
    n1064,
    n913,
    n538,
    n781,
    n384
  );


  xor
  g1128
  (
    n1470,
    n826,
    n886,
    n791,
    n772
  );


  or
  g1129
  (
    n1573,
    n508,
    n499,
    n484,
    n607
  );


  xnor
  g1130
  (
    n1446,
    n769,
    n554,
    n448,
    n524
  );


  and
  g1131
  (
    n1544,
    n824,
    n753,
    n706,
    n606
  );


  xnor
  g1132
  (
    n1550,
    n923,
    n898,
    n513,
    n952
  );


  nand
  g1133
  (
    n1231,
    n883,
    n714,
    n885,
    n874
  );


  nand
  g1134
  (
    n1562,
    n565,
    n566,
    n796,
    n855
  );


  and
  g1135
  (
    n1353,
    n386,
    n779,
    n500,
    n522
  );


  xnor
  g1136
  (
    n1056,
    n675,
    n806,
    n732,
    n494
  );


  xor
  g1137
  (
    n1362,
    n749,
    n925,
    n517,
    n767
  );


  nor
  g1138
  (
    n1401,
    n407,
    n898,
    n394,
    n825
  );


  xnor
  g1139
  (
    n1250,
    n942,
    n473,
    n745,
    n837
  );


  nor
  g1140
  (
    n1390,
    n532,
    n684,
    n487,
    n609
  );


  nor
  g1141
  (
    n1394,
    n550,
    n773,
    n580,
    n395
  );


  nand
  g1142
  (
    n1503,
    n783,
    n895,
    n869,
    n654
  );


  and
  g1143
  (
    n1204,
    n668,
    n708,
    n691,
    n673
  );


  or
  g1144
  (
    n1295,
    n410,
    n448,
    n397,
    n756
  );


  nor
  g1145
  (
    n1106,
    n802,
    n615,
    n449,
    n423
  );


  nor
  g1146
  (
    n1198,
    n544,
    n781,
    n430,
    n401
  );


  nand
  g1147
  (
    n1440,
    n847,
    n575,
    n491,
    n662
  );


  nor
  g1148
  (
    n1546,
    n521,
    n748,
    n910,
    n974
  );


  xnor
  g1149
  (
    n1532,
    n584,
    n763,
    n770,
    n401
  );


  and
  g1150
  (
    n1595,
    n453,
    n961,
    n806,
    n493
  );


  nor
  g1151
  (
    n1148,
    n437,
    n677,
    n830,
    n736
  );


  xor
  g1152
  (
    n1552,
    n573,
    n613,
    n924,
    n499
  );


  xnor
  g1153
  (
    n1115,
    n531,
    n780,
    n478,
    n966
  );


  and
  g1154
  (
    n1019,
    n403,
    n687,
    n854,
    n788
  );


  xor
  g1155
  (
    n1174,
    n812,
    n976,
    n864,
    n741
  );


  xnor
  g1156
  (
    n1489,
    n824,
    n943,
    n960,
    n433
  );


  nand
  g1157
  (
    n1476,
    n851,
    n694,
    n747,
    n811
  );


  and
  g1158
  (
    n1566,
    n905,
    n449,
    n396,
    n454
  );


  xnor
  g1159
  (
    n1091,
    n475,
    n758,
    n553,
    n836
  );


  or
  g1160
  (
    n1015,
    n486,
    n786,
    n954,
    n934
  );


  xor
  g1161
  (
    n1207,
    n921,
    n469,
    n798,
    n952
  );


  nor
  g1162
  (
    n1134,
    n950,
    n678,
    n890,
    n450
  );


  xnor
  g1163
  (
    n1359,
    n892,
    n471,
    n738,
    n782
  );


  xor
  g1164
  (
    n1563,
    n417,
    n777,
    n719,
    n567
  );


  xor
  g1165
  (
    n1445,
    n644,
    n715,
    n447,
    n981
  );


  and
  g1166
  (
    n1582,
    n482,
    n927,
    n506,
    n768
  );


  xor
  g1167
  (
    n1316,
    n935,
    n951,
    n972,
    n665
  );


  xnor
  g1168
  (
    n1026,
    n842,
    n725,
    n800,
    n784
  );


  nand
  g1169
  (
    n1149,
    n701,
    n978,
    n572,
    n891
  );


  or
  g1170
  (
    n1059,
    n426,
    n426,
    n459,
    n733
  );


  and
  g1171
  (
    n1038,
    n611,
    n678,
    n716,
    n563
  );


  nand
  g1172
  (
    n1568,
    n935,
    n758,
    n686,
    n647
  );


  nand
  g1173
  (
    n1114,
    n980,
    n707,
    n545,
    n959
  );


  xor
  g1174
  (
    n1457,
    n815,
    n605,
    n504,
    n853
  );


  nand
  g1175
  (
    n1567,
    n696,
    n538,
    n528,
    n903
  );


  nor
  g1176
  (
    n1146,
    n760,
    n794,
    n480,
    n797
  );


  or
  g1177
  (
    n1041,
    n901,
    n860,
    n525,
    n676
  );


  xnor
  g1178
  (
    n1098,
    n415,
    n705,
    n776,
    n811
  );


  nor
  g1179
  (
    n1039,
    n440,
    n684,
    n718,
    n632
  );


  and
  g1180
  (
    n1239,
    n702,
    n929,
    n944,
    n653
  );


  xor
  g1181
  (
    n1049,
    n930,
    n724,
    n641,
    n977
  );


  nor
  g1182
  (
    n1524,
    n755,
    n948,
    n604,
    n502
  );


  xor
  g1183
  (
    n1235,
    n896,
    n649,
    n651,
    n684
  );


  xnor
  g1184
  (
    n1074,
    n825,
    n424,
    n831,
    n535
  );


  nand
  g1185
  (
    n1346,
    n449,
    n552,
    n955,
    n765
  );


  nand
  g1186
  (
    n1327,
    n780,
    n911,
    n560,
    n644
  );


  nor
  g1187
  (
    n1047,
    n496,
    n982,
    n569,
    n805
  );


  or
  g1188
  (
    n1393,
    n694,
    n388,
    n935,
    n465
  );


  xor
  g1189
  (
    n1406,
    n969,
    n870,
    n655,
    n513
  );


  or
  g1190
  (
    n1051,
    n900,
    n547,
    n960,
    n843
  );


  nand
  g1191
  (
    n1386,
    n772,
    n789,
    n737,
    n865
  );


  or
  g1192
  (
    n1425,
    n874,
    n576,
    n599,
    n469
  );


  xor
  g1193
  (
    n1010,
    n910,
    n427,
    n586,
    n781
  );


  and
  g1194
  (
    n1542,
    n793,
    n451,
    n452,
    n474
  );


  nor
  g1195
  (
    n1430,
    n536,
    n927,
    n420,
    n679
  );


  and
  g1196
  (
    n1061,
    n459,
    n578,
    n759,
    n634
  );


  and
  g1197
  (
    n1408,
    n860,
    n629,
    n900,
    n804
  );


  xnor
  g1198
  (
    n1388,
    n620,
    n754,
    n638,
    n972
  );


  or
  g1199
  (
    n1450,
    n672,
    n923,
    n653,
    n523
  );


  nor
  g1200
  (
    n1269,
    n662,
    n931,
    n404,
    n893
  );


  xor
  g1201
  (
    n1364,
    n698,
    n957,
    n764,
    n603
  );


  xnor
  g1202
  (
    n1375,
    n907,
    n517,
    n693,
    n786
  );


  and
  g1203
  (
    n1246,
    n431,
    n865,
    n659,
    n632
  );


  nor
  g1204
  (
    n1092,
    n975,
    n791,
    n454,
    n582
  );


  and
  g1205
  (
    n1437,
    n959,
    n515,
    n884,
    n988
  );


  nand
  g1206
  (
    n1124,
    n565,
    n531,
    n418,
    n776
  );


  xnor
  g1207
  (
    n1314,
    n858,
    n742,
    n520,
    n702
  );


  nor
  g1208
  (
    n1403,
    n836,
    n444,
    n687,
    n700
  );


  and
  g1209
  (
    n1153,
    n657,
    n947,
    n474,
    n543
  );


  xnor
  g1210
  (
    n1030,
    n478,
    n771,
    n430,
    n901
  );


  xnor
  g1211
  (
    n1287,
    n431,
    n581,
    n472,
    n780
  );


  and
  g1212
  (
    n1116,
    n404,
    n662,
    n717,
    n648
  );


  or
  g1213
  (
    n1385,
    n653,
    n947,
    n907,
    n645
  );


  xnor
  g1214
  (
    n1300,
    n809,
    n712,
    n510,
    n489
  );


  nor
  g1215
  (
    n1119,
    n725,
    n861,
    n583,
    n736
  );


  or
  g1216
  (
    n1551,
    n759,
    n745,
    n550,
    n968
  );


  nand
  g1217
  (
    n1105,
    n559,
    n514,
    n627,
    n843
  );


  xnor
  g1218
  (
    n1182,
    n780,
    n987,
    n949,
    n383
  );


  or
  g1219
  (
    n1065,
    n686,
    n532,
    n828,
    n403
  );


  xor
  g1220
  (
    n1307,
    n966,
    n731,
    n451,
    n967
  );


  nand
  g1221
  (
    n1333,
    n660,
    n701,
    n487,
    n940
  );


  nand
  g1222
  (
    n1428,
    n753,
    n461,
    n882,
    n633
  );


  xnor
  g1223
  (
    n1432,
    n897,
    n694,
    n427,
    n481
  );


  or
  g1224
  (
    n1466,
    n494,
    n751,
    n920,
    n555
  );


  nand
  g1225
  (
    n1495,
    n831,
    n729,
    n871,
    n503
  );


  nor
  g1226
  (
    n1588,
    n538,
    n617,
    n543,
    n561
  );


  xnor
  g1227
  (
    n1221,
    n411,
    n624,
    n925,
    n847
  );


  nand
  g1228
  (
    n1254,
    n625,
    n387,
    n984,
    n533
  );


  xnor
  g1229
  (
    n1277,
    n684,
    n441,
    n890,
    n541
  );


  xor
  g1230
  (
    n1273,
    n623,
    n441,
    n893,
    n795
  );


  nand
  g1231
  (
    n1543,
    n922,
    n876,
    n889,
    n533
  );


  xnor
  g1232
  (
    n1504,
    n469,
    n941,
    n829,
    n872
  );


  xnor
  g1233
  (
    n1130,
    n606,
    n919,
    n570,
    n903
  );


  xor
  g1234
  (
    n1131,
    n400,
    n549,
    n983,
    n847
  );


  xor
  g1235
  (
    n1262,
    n804,
    n630,
    n953,
    n763
  );


  nand
  g1236
  (
    n1426,
    n440,
    n890,
    n900,
    n619
  );


  and
  g1237
  (
    n1554,
    n565,
    n981,
    n954,
    n985
  );


  or
  g1238
  (
    n1444,
    n589,
    n697,
    n728,
    n866
  );


  or
  g1239
  (
    n1058,
    n464,
    n663,
    n575,
    n654
  );


  xnor
  g1240
  (
    n1172,
    n510,
    n731,
    n922,
    n697
  );


  nand
  g1241
  (
    n1150,
    n851,
    n693,
    n911,
    n987
  );


  or
  g1242
  (
    n1305,
    n808,
    n656,
    n432,
    n672
  );


  xnor
  g1243
  (
    n1539,
    n428,
    n518,
    n924,
    n838
  );


  xor
  g1244
  (
    n1145,
    n880,
    n696,
    n399,
    n872
  );


  xnor
  g1245
  (
    n1219,
    n898,
    n635,
    n705,
    n842
  );


  nor
  g1246
  (
    n1270,
    n658,
    n594,
    n568,
    n767
  );


  or
  g1247
  (
    n1226,
    n504,
    n827,
    n475,
    n702
  );


  xor
  g1248
  (
    n1156,
    n846,
    n660,
    n558,
    n937
  );


  nand
  g1249
  (
    n1245,
    n886,
    n595,
    n493,
    n637
  );


  or
  g1250
  (
    n1224,
    n547,
    n921,
    n697,
    n934
  );


  nand
  g1251
  (
    n1220,
    n638,
    n748,
    n857,
    n473
  );


  or
  g1252
  (
    n1215,
    n636,
    n824,
    n915,
    n630
  );


  nor
  g1253
  (
    n1308,
    n645,
    n756,
    n896,
    n738
  );


  and
  g1254
  (
    n1518,
    n432,
    n961,
    n944,
    n654
  );


  or
  g1255
  (
    n1421,
    n627,
    n836,
    n501,
    n690
  );


  and
  g1256
  (
    n1126,
    n988,
    n827,
    n590,
    n595
  );


  or
  g1257
  (
    n1586,
    n952,
    n835,
    n825,
    n600
  );


  xor
  g1258
  (
    n1228,
    n747,
    n908,
    n477,
    n815
  );


  xnor
  g1259
  (
    n1526,
    n785,
    n681,
    n616,
    n751
  );


  nand
  g1260
  (
    n1443,
    n926,
    n940,
    n439,
    n528
  );


  nand
  g1261
  (
    n1397,
    n739,
    n592,
    n486,
    n771
  );


  or
  g1262
  (
    n1487,
    n842,
    n944,
    n679,
    n712
  );


  nor
  g1263
  (
    n1101,
    n574,
    n741,
    n683,
    n965
  );


  and
  g1264
  (
    n1427,
    n689,
    n467,
    n483,
    n949
  );


  xor
  g1265
  (
    n1206,
    n575,
    n546,
    n741,
    n457
  );


  and
  g1266
  (
    n1044,
    n566,
    n669,
    n818,
    n422
  );


  or
  g1267
  (
    n1078,
    n869,
    n614,
    n516,
    n593
  );


  xnor
  g1268
  (
    n1335,
    n450,
    n537,
    n875,
    n906
  );


  xnor
  g1269
  (
    n1311,
    n902,
    n590,
    n557,
    n769
  );


  xor
  g1270
  (
    n1285,
    n748,
    n699,
    n866,
    n884
  );


  nor
  g1271
  (
    n1508,
    n794,
    n507,
    n400,
    n729
  );


  nand
  g1272
  (
    n1136,
    n912,
    n615,
    n513,
    n584
  );


  and
  g1273
  (
    n1138,
    n968,
    n480,
    n622,
    n788
  );


  nor
  g1274
  (
    n1348,
    n820,
    n852,
    n640,
    n730
  );


  nor
  g1275
  (
    n1460,
    n906,
    n586,
    n687,
    n769
  );


  xor
  g1276
  (
    n1334,
    n438,
    n435,
    n785,
    n757
  );


  and
  g1277
  (
    n1167,
    n555,
    n936,
    n779,
    n610
  );


  nand
  g1278
  (
    n1459,
    n746,
    n786,
    n583,
    n674
  );


  or
  g1279
  (
    n1547,
    n816,
    n571,
    n464,
    n428
  );


  nor
  g1280
  (
    n1448,
    n576,
    n887,
    n706,
    n489
  );


  xnor
  g1281
  (
    n1248,
    n871,
    n564,
    n601,
    n807
  );


  or
  g1282
  (
    n1493,
    n440,
    n652,
    n877,
    n497
  );


  or
  g1283
  (
    n1572,
    n678,
    n802,
    n881,
    n899
  );


  or
  g1284
  (
    n1431,
    n650,
    n832,
    n614,
    n948
  );


  nand
  g1285
  (
    n1356,
    n978,
    n470,
    n957,
    n373
  );


  nand
  g1286
  (
    n1447,
    n668,
    n955,
    n481,
    n861
  );


  nor
  g1287
  (
    n1183,
    n580,
    n377,
    n651,
    n490
  );


  or
  g1288
  (
    n1441,
    n485,
    n856,
    n699,
    n521
  );


  nand
  g1289
  (
    n1280,
    n919,
    n710,
    n436,
    n665
  );


  nand
  g1290
  (
    n1400,
    n589,
    n525,
    n501,
    n421
  );


  xnor
  g1291
  (
    n1293,
    n525,
    n690,
    n945,
    n755
  );


  or
  g1292
  (
    n1147,
    n886,
    n600,
    n782,
    n633
  );


  and
  g1293
  (
    n1094,
    n754,
    n709,
    n510,
    n908
  );


  nor
  g1294
  (
    n1166,
    n971,
    n645,
    n509,
    n893
  );


  nor
  g1295
  (
    n1347,
    n616,
    n949,
    n548,
    n471
  );


  xnor
  g1296
  (
    n1350,
    n917,
    n880,
    n963,
    n581
  );


  nor
  g1297
  (
    n1029,
    n596,
    n784,
    n722,
    n793
  );


  xnor
  g1298
  (
    n1374,
    n840,
    n962,
    n580,
    n971
  );


  or
  g1299
  (
    n1195,
    n634,
    n463,
    n937,
    n984
  );


  xnor
  g1300
  (
    n1046,
    n670,
    n881,
    n927,
    n838
  );


  or
  g1301
  (
    n1160,
    n412,
    n602,
    n604,
    n798
  );


  or
  g1302
  (
    n1276,
    n873,
    n616,
    n502,
    n743
  );


  nand
  g1303
  (
    n1391,
    n477,
    n764,
    n636,
    n904
  );


  or
  g1304
  (
    n1575,
    n721,
    n963,
    n599,
    n505
  );


  xnor
  g1305
  (
    n1034,
    n573,
    n942,
    n704,
    n922
  );


  and
  g1306
  (
    n1358,
    n438,
    n968,
    n475,
    n986
  );


  and
  g1307
  (
    n1462,
    n658,
    n399,
    n442,
    n588
  );


  nor
  g1308
  (
    n1414,
    n916,
    n688,
    n856,
    n734
  );


  xor
  g1309
  (
    n1159,
    n611,
    n728,
    n540,
    n787
  );


  nor
  g1310
  (
    n1468,
    n655,
    n974,
    n525,
    n833
  );


  nor
  g1311
  (
    n1144,
    n658,
    n962,
    n898,
    n696
  );


  and
  g1312
  (
    n1389,
    n559,
    n819,
    n579,
    n946
  );


  nand
  g1313
  (
    n1143,
    n514,
    n866,
    n805,
    n678
  );


  and
  g1314
  (
    n1553,
    n546,
    n688,
    n519,
    n518
  );


  xnor
  g1315
  (
    n1520,
    n969,
    n777,
    n844,
    n911
  );


  xnor
  g1316
  (
    n1178,
    n829,
    n916,
    n443,
    n848
  );


  or
  g1317
  (
    n1112,
    n826,
    n499,
    n935,
    n586
  );


  xnor
  g1318
  (
    n1332,
    n513,
    n897,
    n909,
    n621
  );


  or
  g1319
  (
    n1188,
    n500,
    n516,
    n961,
    n428
  );


  nand
  g1320
  (
    n1383,
    n393,
    n926,
    n883,
    n807
  );


  xnor
  g1321
  (
    n1294,
    n650,
    n565,
    n456,
    n558
  );


  nand
  g1322
  (
    n1324,
    n647,
    n980,
    n412,
    n520
  );


  nor
  g1323
  (
    n1505,
    n853,
    n919,
    n498,
    n752
  );


  xor
  g1324
  (
    n1090,
    n951,
    n735,
    n622,
    n520
  );


  or
  g1325
  (
    n1410,
    n705,
    n938,
    n917,
    n597
  );


  xnor
  g1326
  (
    n1339,
    n824,
    n745,
    n437,
    n481
  );


  nor
  g1327
  (
    n1472,
    n790,
    n757,
    n792,
    n443
  );


  xor
  g1328
  (
    n1129,
    n568,
    n682,
    n877,
    n943
  );


  or
  g1329
  (
    n1066,
    n603,
    n579,
    n723,
    n424
  );


  xnor
  g1330
  (
    n1125,
    n681,
    n915,
    n818,
    n876
  );


  nor
  g1331
  (
    n1590,
    n398,
    n883,
    n605,
    n856
  );


  xnor
  g1332
  (
    n1453,
    n912,
    n447,
    n472,
    n749
  );


  nand
  g1333
  (
    n1249,
    n877,
    n504,
    n539,
    n816
  );


  nor
  g1334
  (
    n1140,
    n574,
    n712,
    n560,
    n463
  );


  nand
  g1335
  (
    n1292,
    n871,
    n703,
    n566,
    n577
  );


  or
  g1336
  (
    n1108,
    n467,
    n834,
    n956,
    n414
  );


  nand
  g1337
  (
    n1558,
    n644,
    n926,
    n663,
    n919
  );


  xor
  g1338
  (
    n1263,
    n723,
    n924,
    n892,
    n578
  );


  nor
  g1339
  (
    n1405,
    n474,
    n659,
    n465,
    n903
  );


  or
  g1340
  (
    n1110,
    n804,
    n708,
    n974,
    n495
  );


  nand
  g1341
  (
    n1152,
    n605,
    n914,
    n827,
    n492
  );


  xor
  g1342
  (
    n1286,
    n464,
    n534,
    n689,
    n693
  );


  xnor
  g1343
  (
    n1012,
    n675,
    n876,
    n420,
    n544
  );


  xor
  g1344
  (
    n1564,
    n809,
    n734,
    n526,
    n585
  );


  nand
  g1345
  (
    n1222,
    n854,
    n372,
    n931,
    n646
  );


  and
  g1346
  (
    n1591,
    n718,
    n767,
    n594,
    n836
  );


  and
  g1347
  (
    n1415,
    n673,
    n759,
    n382,
    n868
  );


  xnor
  g1348
  (
    n1100,
    n891,
    n685,
    n768,
    n985
  );


  or
  g1349
  (
    n1244,
    n381,
    n729,
    n977,
    n742
  );


  xor
  g1350
  (
    n1075,
    n529,
    n496,
    n488,
    n713
  );


  xor
  g1351
  (
    n1265,
    n764,
    n844,
    n472,
    n531
  );


  nand
  g1352
  (
    n1517,
    n868,
    n666,
    n755,
    n806
  );


  or
  g1353
  (
    n1168,
    n810,
    n885,
    n636,
    n930
  );


  xnor
  g1354
  (
    n1072,
    n466,
    n869,
    n691,
    n835
  );


  xnor
  g1355
  (
    n1545,
    n867,
    n609,
    n641,
    n785
  );


  or
  g1356
  (
    n1531,
    n846,
    n792,
    n834,
    n704
  );


  nor
  g1357
  (
    n1514,
    n445,
    n453,
    n925,
    n483
  );


  xor
  g1358
  (
    n1021,
    n817,
    n434,
    n458,
    n733
  );


  and
  g1359
  (
    n1133,
    n940,
    n975,
    n637,
    n526
  );


  nand
  g1360
  (
    n1201,
    n970,
    n965,
    n429,
    n911
  );


  xnor
  g1361
  (
    n1256,
    n710,
    n452,
    n778,
    n833
  );


  and
  g1362
  (
    n1373,
    n680,
    n641,
    n660,
    n844
  );


  xor
  g1363
  (
    n1519,
    n710,
    n424,
    n843,
    n518
  );


  xor
  g1364
  (
    n1020,
    n436,
    n717,
    n497,
    n468
  );


  nor
  g1365
  (
    n1474,
    n873,
    n650,
    n571,
    n762
  );


  xnor
  g1366
  (
    n1378,
    n505,
    n577,
    n872,
    n916
  );


  nand
  g1367
  (
    n1337,
    n858,
    n665,
    n769,
    n771
  );


  xor
  g1368
  (
    n1309,
    n631,
    n495,
    n751,
    n832
  );


  nand
  g1369
  (
    n1236,
    n899,
    n831,
    n497,
    n402
  );


  or
  g1370
  (
    n1118,
    n530,
    n839,
    n611,
    n867
  );


  and
  g1371
  (
    n1392,
    n956,
    n749,
    n533,
    n407
  );


  nand
  g1372
  (
    n1483,
    n691,
    n425,
    n985,
    n557
  );


  nand
  g1373
  (
    n1216,
    n535,
    n976,
    n631,
    n861
  );


  and
  g1374
  (
    n1371,
    n567,
    n725,
    n944,
    n679
  );


  nor
  g1375
  (
    n1541,
    n671,
    n988,
    n623,
    n527
  );


  xor
  g1376
  (
    n1103,
    n813,
    n456,
    n731,
    n907
  );


  or
  g1377
  (
    n1243,
    n673,
    n619,
    n796,
    n621
  );


  nand
  g1378
  (
    n1128,
    n967,
    n550,
    n460,
    n472
  );


  xnor
  g1379
  (
    n1433,
    n728,
    n683,
    n406,
    n815
  );


  nand
  g1380
  (
    n1199,
    n948,
    n556,
    n821,
    n598
  );


  nor
  g1381
  (
    n1491,
    n742,
    n852,
    n914,
    n768
  );


  or
  g1382
  (
    n1369,
    n984,
    n772,
    n553,
    n508
  );


  nor
  g1383
  (
    n1192,
    n389,
    n446,
    n888,
    n760
  );


  xor
  g1384
  (
    n1027,
    n841,
    n908,
    n508,
    n948
  );


  nor
  g1385
  (
    n1571,
    n608,
    n433,
    n711,
    n612
  );


  xor
  g1386
  (
    n1434,
    n889,
    n930,
    n545,
    n981
  );


  nor
  g1387
  (
    n1429,
    n887,
    n425,
    n496,
    n482
  );


  nor
  g1388
  (
    n1565,
    n777,
    n641,
    n692,
    n863
  );


  or
  g1389
  (
    n1296,
    n546,
    n889,
    n857,
    n485
  );


  xnor
  g1390
  (
    n1458,
    n564,
    n462,
    n743,
    n544
  );


  and
  g1391
  (
    n1083,
    n475,
    n833,
    n502,
    n501
  );


  xor
  g1392
  (
    n1151,
    n859,
    n908,
    n803,
    n989
  );


  xnor
  g1393
  (
    n1288,
    n547,
    n697,
    n651,
    n628
  );


  xor
  g1394
  (
    n1502,
    n867,
    n708,
    n934,
    n647
  );


  xnor
  g1395
  (
    n1328,
    n726,
    n514,
    n536,
    n762
  );


  xnor
  g1396
  (
    n1379,
    n737,
    n928,
    n868,
    n650
  );


  xor
  g1397
  (
    n1321,
    n443,
    n686,
    n803,
    n761
  );


  xor
  g1398
  (
    n1086,
    n492,
    n438,
    n713,
    n495
  );


  nand
  g1399
  (
    n1329,
    n587,
    n501,
    n671,
    n466
  );


  nor
  g1400
  (
    n1281,
    n720,
    n978,
    n647,
    n657
  );


  or
  g1401
  (
    n1326,
    n839,
    n736,
    n593,
    n459
  );


  nand
  g1402
  (
    n1197,
    n928,
    n884,
    n762,
    n894
  );


  or
  g1403
  (
    n1454,
    n512,
    n978,
    n976,
    n964
  );


  xor
  g1404
  (
    n1578,
    n765,
    n823,
    n676,
    n804
  );


  nand
  g1405
  (
    n1011,
    n829,
    n913,
    n429,
    n431
  );


  xor
  g1406
  (
    n1202,
    n558,
    n802,
    n958,
    n709
  );


  xnor
  g1407
  (
    n1384,
    n687,
    n941,
    n595,
    n761
  );


  nand
  g1408
  (
    n1576,
    n820,
    n987,
    n691,
    n743
  );


  and
  g1409
  (
    n1496,
    n733,
    n826,
    n524,
    n626
  );


  xnor
  g1410
  (
    n1259,
    n901,
    n891,
    n442,
    n619
  );


  xor
  g1411
  (
    n1506,
    n771,
    n667,
    n762,
    n433
  );


  nor
  g1412
  (
    n1511,
    n725,
    n910,
    n881,
    n863
  );


  and
  g1413
  (
    n1205,
    n452,
    n801,
    n593,
    n904
  );


  nor
  g1414
  (
    n1171,
    n628,
    n675,
    n535,
    n797
  );


  and
  g1415
  (
    n1480,
    n879,
    n538,
    n622,
    n503
  );


  nand
  g1416
  (
    n1331,
    n556,
    n588,
    n484,
    n975
  );


  xnor
  g1417
  (
    n1407,
    n524,
    n889,
    n598,
    n632
  );


  or
  g1418
  (
    n1229,
    n503,
    n448,
    n875,
    n649
  );


  xnor
  g1419
  (
    n1196,
    n628,
    n685,
    n529,
    n930
  );


  nand
  g1420
  (
    n1510,
    n572,
    n921,
    n480,
    n548
  );


  nor
  g1421
  (
    n1561,
    n744,
    n534,
    n460,
    n698
  );


  and
  g1422
  (
    n1577,
    n832,
    n458,
    n419,
    n801
  );


  and
  g1423
  (
    n1357,
    n441,
    n834,
    n953,
    n591
  );


  nor
  g1424
  (
    n1592,
    n857,
    n568,
    n552,
    n880
  );


  nand
  g1425
  (
    n1525,
    n610,
    n559,
    n530,
    n444
  );


  nand
  g1426
  (
    n1088,
    n643,
    n673,
    n542,
    n979
  );


  xnor
  g1427
  (
    n1186,
    n939,
    n914,
    n853,
    n664
  );


  nand
  g1428
  (
    n1233,
    n576,
    n665,
    n808,
    n850
  );


  nor
  g1429
  (
    n1319,
    n643,
    n796,
    n380,
    n983
  );


  xnor
  g1430
  (
    n1419,
    n698,
    n949,
    n447,
    n479
  );


  nand
  g1431
  (
    n1313,
    n704,
    n776,
    n522,
    n819
  );


  nor
  g1432
  (
    n1063,
    n634,
    n808,
    n554,
    n779
  );


  and
  g1433
  (
    n1014,
    n635,
    n457,
    n878,
    n705
  );


  xor
  g1434
  (
    n1025,
    n695,
    n778,
    n957,
    n816
  );


  xnor
  g1435
  (
    n1102,
    n670,
    n439,
    n539
  );


  xnor
  g1436
  (
    n1521,
    n854,
    n761,
    n983,
    n708
  );


  or
  g1437
  (
    n1241,
    n833,
    n852,
    n962,
    n927
  );


  nor
  g1438
  (
    n1536,
    n901,
    n692,
    n800,
    n966
  );


  xnor
  g1439
  (
    n1037,
    n941,
    n936,
    n925,
    n822
  );


  xnor
  g1440
  (
    n1549,
    n408,
    n845,
    n655,
    n616
  );


  and
  g1441
  (
    n1022,
    n508,
    n763,
    n795,
    n951
  );


  and
  g1442
  (
    n1104,
    n654,
    n962,
    n937,
    n707
  );


  or
  g1443
  (
    n1121,
    n635,
    n682,
    n505,
    n895
  );


  nor
  g1444
  (
    n1067,
    n445,
    n711,
    n863,
    n768
  );


  xor
  g1445
  (
    n1055,
    n466,
    n540,
    n872,
    n630
  );


  xnor
  g1446
  (
    n1485,
    n573,
    n933,
    n530,
    n690
  );


  and
  g1447
  (
    n1267,
    n664,
    n456,
    n740,
    n482
  );


  or
  g1448
  (
    n1409,
    n862,
    n707,
    n427,
    n523
  );


  xnor
  g1449
  (
    n1312,
    n587,
    n766,
    n852,
    n557
  );


  xnor
  g1450
  (
    n1289,
    n488,
    n413,
    n955,
    n569
  );


  or
  g1451
  (
    n1238,
    n434,
    n938,
    n455,
    n813
  );


  and
  g1452
  (
    n1070,
    n563,
    n724,
    n527,
    n799
  );


  nand
  g1453
  (
    n1497,
    n648,
    n507,
    n840,
    n542
  );


  xor
  g1454
  (
    n1560,
    n865,
    n942,
    n455,
    n757
  );


  xnor
  g1455
  (
    n1208,
    n506,
    n793,
    n895,
    n590
  );


  and
  g1456
  (
    n1031,
    n623,
    n828,
    n848,
    n774
  );


  or
  g1457
  (
    n1360,
    n603,
    n637,
    n445,
    n965
  );


  nand
  g1458
  (
    n1507,
    n479,
    n617,
    n459,
    n474
  );


  xor
  g1459
  (
    n1099,
    n455,
    n683,
    n620,
    n625
  );


  and
  g1460
  (
    n1062,
    n722,
    n989,
    n888,
    n937
  );


  nor
  g1461
  (
    n1317,
    n720,
    n649,
    n730,
    n727
  );


  nand
  g1462
  (
    n1093,
    n913,
    n873,
    n700,
    n932
  );


  and
  g1463
  (
    n1290,
    n721,
    n528,
    n958,
    n947
  );


  nand
  g1464
  (
    n1085,
    n628,
    n462,
    n391,
    n734
  );


  nand
  g1465
  (
    n1352,
    n376,
    n808,
    n671,
    n969
  );


  nor
  g1466
  (
    n1424,
    n589,
    n408,
    n820,
    n870
  );


  nand
  g1467
  (
    n1271,
    n435,
    n738,
    n835,
    n629
  );


  xor
  g1468
  (
    n1173,
    n505,
    n449,
    n798,
    n543
  );


  nand
  g1469
  (
    n1185,
    n522,
    n591,
    n421,
    n531
  );


  nand
  g1470
  (
    n1218,
    n770,
    n473,
    n756,
    n583
  );


  nand
  g1471
  (
    n1096,
    n468,
    n713,
    n773,
    n740
  );


  nand
  g1472
  (
    n1180,
    n588,
    n405,
    n506,
    n810
  );


  xnor
  g1473
  (
    n1252,
    n669,
    n447,
    n544,
    n592
  );


  and
  g1474
  (
    n1323,
    n928,
    n629,
    n506,
    n760
  );


  nand
  g1475
  (
    n1585,
    n642,
    n853,
    n818,
    n556
  );


  or
  g1476
  (
    n1482,
    n692,
    n918,
    n637,
    n509
  );


  and
  g1477
  (
    n1177,
    n721,
    n875,
    n640,
    n570
  );


  nand
  g1478
  (
    n1053,
    n781,
    n518,
    n596,
    n434
  );


  xor
  g1479
  (
    n1529,
    n846,
    n390,
    n648,
    n444
  );


  nand
  g1480
  (
    n1556,
    n823,
    n488,
    n612,
    n371
  );


  nor
  g1481
  (
    n1417,
    n638,
    n580,
    n718,
    n561
  );


  or
  g1482
  (
    n1367,
    n913,
    n446,
    n891,
    n490
  );


  nand
  g1483
  (
    n1117,
    n436,
    n902,
    n527,
    n483
  );


  xnor
  g1484
  (
    n1442,
    n977,
    n416,
    n601,
    n589
  );


  nand
  g1485
  (
    n1165,
    n677,
    n942,
    n701,
    n375
  );


  xor
  g1486
  (
    n1033,
    n572,
    n601,
    n667,
    n584
  );


  nand
  g1487
  (
    n1135,
    n631,
    n555,
    n618,
    n960
  );


  or
  g1488
  (
    n1381,
    n389,
    n468,
    n618,
    n834
  );


  xnor
  g1489
  (
    n1122,
    n643,
    n562,
    n488,
    n775
  );


  nor
  g1490
  (
    n1068,
    n614,
    n651,
    n549,
    n841
  );


  or
  g1491
  (
    n1097,
    n624,
    n774,
    n915,
    n945
  );


  and
  g1492
  (
    n1212,
    n668,
    n570,
    n619,
    n838
  );


  nor
  g1493
  (
    n1548,
    n830,
    n548,
    n682,
    n639
  );


  and
  g1494
  (
    n1435,
    n805,
    n466,
    n642,
    n553
  );


  xor
  g1495
  (
    n1523,
    n435,
    n786,
    n652,
    n693
  );


  and
  g1496
  (
    n1372,
    n814,
    n515,
    n787,
    n761
  );


  xnor
  g1497
  (
    n1282,
    n982,
    n405,
    n918,
    n618
  );


  xor
  g1498
  (
    n1478,
    n720,
    n918,
    n500,
    n867
  );


  xor
  g1499
  (
    n1593,
    n736,
    n918,
    n549,
    n764
  );


  or
  g1500
  (
    n1298,
    n566,
    n624,
    n585,
    n887
  );


  or
  g1501
  (
    n1513,
    n666,
    n511,
    n929,
    n951
  );


  or
  g1502
  (
    n1230,
    n395,
    n814,
    n575,
    n907
  );


  and
  g1503
  (
    n1533,
    n451,
    n738,
    n504,
    n397
  );


  or
  g1504
  (
    n1574,
    n952,
    n409,
    n625,
    n695
  );


  and
  g1505
  (
    n1528,
    n479,
    n577,
    n631,
    n848
  );


  nor
  g1506
  (
    n1481,
    n939,
    n478,
    n849,
    n984
  );


  nor
  g1507
  (
    n1162,
    n954,
    n839,
    n947,
    n921
  );


  or
  g1508
  (
    n1194,
    n767,
    n563,
    n766,
    n752
  );


  xnor
  g1509
  (
    n1535,
    n591,
    n646,
    n939,
    n672
  );


  and
  g1510
  (
    n1123,
    n874,
    n788,
    n960,
    n498
  );


  or
  g1511
  (
    n1191,
    n815,
    n963,
    n932,
    n510
  );


  and
  g1512
  (
    n1132,
    n677,
    n760,
    n599,
    n515
  );


  xnor
  g1513
  (
    n1213,
    n838,
    n706,
    n979,
    n874
  );


  nor
  g1514
  (
    n1193,
    n646,
    n652,
    n436,
    n648
  );


  nand
  g1515
  (
    n1423,
    n756,
    n613,
    n865,
    n423
  );


  xor
  g1516
  (
    n1043,
    n432,
    n883,
    n822,
    n970
  );


  xnor
  g1517
  (
    n1109,
    n441,
    n676,
    n791,
    n847
  );


  nand
  g1518
  (
    n1073,
    n744,
    n470,
    n976,
    n809
  );


  nand
  g1519
  (
    n1322,
    n724,
    n653,
    n854,
    n775
  );


  nor
  g1520
  (
    n1057,
    n439,
    n982,
    n763,
    n430
  );


  or
  g1521
  (
    n1175,
    n703,
    n807,
    n463,
    n811
  );


  nand
  g1522
  (
    n1420,
    n489,
    n529,
    n851,
    n670
  );


  nor
  g1523
  (
    n1141,
    n512,
    n617,
    n972,
    n726
  );


  nand
  g1524
  (
    n1155,
    n523,
    n542,
    n827,
    n766
  );


  or
  g1525
  (
    n1515,
    n892,
    n640,
    n433,
    n986
  );


  xor
  g1526
  (
    n1258,
    n792,
    n541,
    n888,
    n604
  );


  xor
  g1527
  (
    n1275,
    n495,
    n926,
    n723,
    n953
  );


  xnor
  g1528
  (
    n1402,
    n849,
    n484,
    n783,
    n774
  );


  xor
  g1529
  (
    n1368,
    n709,
    n929,
    n735,
    n750
  );


  xor
  g1530
  (
    n1268,
    n881,
    n555,
    n602,
    n868
  );


  xor
  g1531
  (
    n1418,
    n524,
    n390,
    n694,
    n884
  );


  xor
  g1532
  (
    n1449,
    n406,
    n778,
    n856,
    n906
  );


  xnor
  g1533
  (
    n1283,
    n920,
    n493,
    n850,
    n812
  );


  nor
  g1534
  (
    n1594,
    n864,
    n370,
    n568,
    n974
  );


  xnor
  g1535
  (
    n1455,
    n902,
    n511,
    n526,
    n882
  );


  nor
  g1536
  (
    n1471,
    n458,
    n583,
    n640,
    n800
  );


  xor
  g1537
  (
    n1343,
    n630,
    n957,
    n845,
    n732
  );


  nand
  g1538
  (
    n1349,
    n460,
    n457,
    n817,
    n627
  );


  xor
  g1539
  (
    n1018,
    n879,
    n924,
    n587,
    n462
  );


  xor
  g1540
  (
    n1050,
    n674,
    n787,
    n840,
    n803
  );


  nand
  g1541
  (
    n1107,
    n855,
    n714,
    n558,
    n765
  );


  and
  g1542
  (
    n1579,
    n391,
    n541,
    n668,
    n923
  );


  nand
  g1543
  (
    n1538,
    n701,
    n775,
    n610,
    n446
  );


  xor
  g1544
  (
    n1016,
    n590,
    n970,
    n715,
    n576
  );


  xnor
  g1545
  (
    n1161,
    n644,
    n663,
    n794,
    n517
  );


  nand
  g1546
  (
    n1080,
    n489,
    n465,
    n659,
    n740
  );


  xor
  g1547
  (
    n1036,
    n928,
    n543,
    n846,
    n470
  );


  and
  g1548
  (
    n1013,
    n607,
    n666,
    n633,
    n396
  );


  xor
  g1549
  (
    n1501,
    n638,
    n801,
    n582,
    n826
  );


  xnor
  g1550
  (
    n1411,
    n415,
    n432,
    n855,
    n430
  );


  or
  g1551
  (
    n1023,
    n912,
    n540,
    n581,
    n841
  );


  nor
  g1552
  (
    n1488,
    n669,
    n699,
    n746,
    n553
  );


  xnor
  g1553
  (
    n1176,
    n551,
    n707,
    n821,
    n969
  );


  nor
  g1554
  (
    n1399,
    n950,
    n388,
    n757,
    n530
  );


  nand
  g1555
  (
    n1082,
    n608,
    n440,
    n909,
    n904
  );


  xnor
  g1556
  (
    n1469,
    n561,
    n737,
    n885,
    n791
  );


  nand
  g1557
  (
    n1232,
    n753,
    n498,
    n567,
    n931
  );


  and
  g1558
  (
    n1247,
    n562,
    n477,
    n626,
    n839
  );


  xnor
  g1559
  (
    n1095,
    n689,
    n799,
    n461,
    n536
  );


  nand
  g1560
  (
    n1297,
    n674,
    n747,
    n759,
    n850
  );


  xor
  g1561
  (
    n1306,
    n548,
    n946,
    n727,
    n858
  );


  nand
  g1562
  (
    n1069,
    n520,
    n680,
    n743,
    n896
  );


  nand
  g1563
  (
    n1475,
    n562,
    n607,
    n821,
    n971
  );


  and
  g1564
  (
    n1341,
    n933,
    n635,
    n784,
    n894
  );


  nor
  g1565
  (
    n1690,
    n1183,
    n1289,
    n1247,
    n1031
  );


  or
  g1566
  (
    n1613,
    n1379,
    n1078,
    n1371,
    n1354
  );


  and
  g1567
  (
    n1646,
    n1036,
    n1053,
    n1037,
    n1215
  );


  or
  g1568
  (
    n1680,
    n1178,
    n1137,
    n1106,
    n1233
  );


  or
  g1569
  (
    n1672,
    n1139,
    n1281,
    n1203,
    n1262
  );


  and
  g1570
  (
    n1640,
    n1389,
    n1111,
    n1388,
    n1227
  );


  nor
  g1571
  (
    n1611,
    n1368,
    n1150,
    n1153,
    n1076
  );


  or
  g1572
  (
    n1676,
    n1017,
    n1392,
    n1278,
    n1243
  );


  nand
  g1573
  (
    n1608,
    n1174,
    n1093,
    n1302,
    n1077
  );


  xnor
  g1574
  (
    n1629,
    n1056,
    n1142,
    n1299,
    n1383
  );


  xnor
  g1575
  (
    n1643,
    n1030,
    n1282,
    n1026,
    n1134
  );


  nand
  g1576
  (
    n1678,
    n1016,
    n1200,
    n1387,
    n1068
  );


  nand
  g1577
  (
    n1691,
    n1204,
    n1167,
    n1349,
    n1259
  );


  nor
  g1578
  (
    n1674,
    n1164,
    n1390,
    n1171,
    n1350
  );


  or
  g1579
  (
    n1651,
    n1103,
    n1105,
    n1058,
    n1293
  );


  nand
  g1580
  (
    n1644,
    n1019,
    n1273,
    n1249,
    n1198
  );


  and
  g1581
  (
    n1626,
    n1193,
    n1225,
    n1059,
    n1045
  );


  and
  g1582
  (
    n1654,
    n1328,
    n1157,
    n1028,
    n1307
  );


  and
  g1583
  (
    n1658,
    n1329,
    n1377,
    n1009,
    n1197
  );


  xnor
  g1584
  (
    n1624,
    n1086,
    n1365,
    n1100,
    n1035
  );


  xor
  g1585
  (
    n1604,
    n1049,
    n1340,
    n1291,
    n1122
  );


  or
  g1586
  (
    n1609,
    n1163,
    n1113,
    n1337,
    n1060
  );


  or
  g1587
  (
    n1642,
    n1364,
    n1222,
    n1376,
    n1219
  );


  and
  g1588
  (
    n1659,
    n1187,
    n1265,
    n1136,
    n1224
  );


  nor
  g1589
  (
    n1621,
    n1155,
    n1303,
    n1320,
    n1083
  );


  xnor
  g1590
  (
    n1614,
    n1319,
    n1207,
    n1236,
    n1335
  );


  xor
  g1591
  (
    n1683,
    n1088,
    n1089,
    n1324,
    n1067
  );


  and
  g1592
  (
    n1601,
    n1358,
    n1300,
    n1280,
    n1109
  );


  and
  g1593
  (
    n1634,
    n1374,
    n1112,
    n1326,
    n1250
  );


  nand
  g1594
  (
    n1655,
    n1196,
    n1271,
    n1199,
    n1384
  );


  nand
  g1595
  (
    n1664,
    n1101,
    n1373,
    n1217,
    n1190
  );


  nor
  g1596
  (
    n1652,
    n1336,
    n1380,
    n1073,
    n1143
  );


  xnor
  g1597
  (
    n1679,
    n1108,
    n1301,
    n1242,
    n1294
  );


  xnor
  g1598
  (
    n1682,
    n1127,
    n1075,
    n1356,
    n1180
  );


  or
  g1599
  (
    n1662,
    n1375,
    n1235,
    n1051,
    n1208
  );


  and
  g1600
  (
    n1689,
    n1191,
    n1268,
    n1149,
    n1098
  );


  xor
  g1601
  (
    n1623,
    n1241,
    n1325,
    n1161,
    n1274
  );


  xnor
  g1602
  (
    n1630,
    n1091,
    n1168,
    n1085,
    n1355
  );


  and
  g1603
  (
    n1650,
    n1061,
    n1159,
    n1186,
    n1285
  );


  nand
  g1604
  (
    n1599,
    n1033,
    n1366,
    n1270,
    n1170
  );


  xnor
  g1605
  (
    n1632,
    n1039,
    n1216,
    n1211,
    n1116
  );


  nor
  g1606
  (
    n1622,
    n1173,
    n1042,
    n1266,
    n1162
  );


  or
  g1607
  (
    n1692,
    n1359,
    n1027,
    n1125,
    n1040
  );


  nor
  g1608
  (
    n1615,
    n1367,
    n1263,
    n1237,
    n1297
  );


  xor
  g1609
  (
    n1661,
    n1378,
    n1117,
    n1258,
    n1015
  );


  nand
  g1610
  (
    n1617,
    n1070,
    n1012,
    n1124,
    n1129
  );


  or
  g1611
  (
    n1631,
    n1251,
    n1338,
    n1209,
    n1323
  );


  nor
  g1612
  (
    n1668,
    n1231,
    n1057,
    n1210,
    n1309
  );


  and
  g1613
  (
    n1602,
    n1072,
    n1346,
    n1385,
    n1310
  );


  xor
  g1614
  (
    n1648,
    n1052,
    n1110,
    n1321,
    n1351
  );


  xor
  g1615
  (
    n1636,
    n1244,
    n1382,
    n1022,
    n1194
  );


  and
  g1616
  (
    n1620,
    n1032,
    n1014,
    n1316,
    n1331
  );


  xnor
  g1617
  (
    n1645,
    n1205,
    n1314,
    n1094,
    n1317
  );


  or
  g1618
  (
    n1656,
    n1361,
    n1295,
    n1119,
    n1050
  );


  xor
  g1619
  (
    n1637,
    n1283,
    n1029,
    n1107,
    n1195
  );


  xor
  g1620
  (
    n1639,
    n1213,
    n1055,
    n1046,
    n1230
  );


  nor
  g1621
  (
    n1663,
    n1018,
    n1189,
    n1372,
    n1287
  );


  and
  g1622
  (
    n1666,
    n1165,
    n1130,
    n1234,
    n1158
  );


  nor
  g1623
  (
    n1675,
    n1315,
    n1151,
    n1141,
    n1047
  );


  or
  g1624
  (
    n1660,
    n1144,
    n1145,
    n1353,
    n1362
  );


  xor
  g1625
  (
    n1627,
    n1146,
    n1148,
    n1041,
    n1201
  );


  nor
  g1626
  (
    n1677,
    n1298,
    n1126,
    n1175,
    n1084
  );


  xor
  g1627
  (
    n1673,
    n1256,
    n1154,
    n1074,
    n1169
  );


  or
  g1628
  (
    n1618,
    n1232,
    n1104,
    n1275,
    n1087
  );


  and
  g1629
  (
    n1635,
    n1330,
    n1188,
    n1218,
    n1223
  );


  nand
  g1630
  (
    n1606,
    n1080,
    n1357,
    n1363,
    n1184
  );


  and
  g1631
  (
    n1671,
    n1021,
    n1252,
    n1185,
    n1177
  );


  nor
  g1632
  (
    n1628,
    n1115,
    n1114,
    n1081,
    n1128
  );


  nand
  g1633
  (
    n1647,
    n1131,
    n1034,
    n1011,
    n1343
  );


  xor
  g1634
  (
    n1605,
    n1332,
    n1286,
    n1352,
    n1311
  );


  xor
  g1635
  (
    n1641,
    n1288,
    n1024,
    n1069,
    n1092
  );


  nand
  g1636
  (
    n1688,
    n1248,
    n1097,
    n1135,
    n1214
  );


  and
  g1637
  (
    n1616,
    n1239,
    n1176,
    n1202,
    n1381
  );


  nand
  g1638
  (
    n1649,
    n1221,
    n1339,
    n1043,
    n1220
  );


  nor
  g1639
  (
    n1687,
    n1020,
    n1240,
    n1095,
    n1305
  );


  and
  g1640
  (
    n1607,
    n1226,
    n1123,
    n1391,
    n1133
  );


  xnor
  g1641
  (
    n1653,
    n1308,
    n1347,
    n1269,
    n1360
  );


  and
  g1642
  (
    n1633,
    n1260,
    n1192,
    n1264,
    n1296
  );


  nor
  g1643
  (
    n1686,
    n1044,
    n1238,
    n1140,
    n1386
  );


  nand
  g1644
  (
    n1600,
    n1277,
    n1279,
    n1245,
    n1054
  );


  or
  g1645
  (
    n1610,
    n1284,
    n1182,
    n1071,
    n1345
  );


  and
  g1646
  (
    n1638,
    n1065,
    n1096,
    n1257,
    n1267
  );


  or
  g1647
  (
    n1657,
    n1079,
    n1160,
    n1253,
    n1102
  );


  or
  g1648
  (
    n1669,
    n1181,
    n1010,
    n1327,
    n1254
  );


  nand
  g1649
  (
    n1612,
    n1013,
    n1156,
    n1048,
    n1062
  );


  xnor
  g1650
  (
    n1685,
    n1292,
    n1246,
    n1138,
    n1172
  );


  xnor
  g1651
  (
    n1598,
    n1348,
    n1063,
    n1304,
    n1152
  );


  nand
  g1652
  (
    n1619,
    n1333,
    n1025,
    n1306,
    n1228
  );


  nand
  g1653
  (
    n1665,
    n1121,
    n1118,
    n1147,
    n1206
  );


  xor
  g1654
  (
    n1603,
    n1082,
    n1369,
    n1272,
    n1064
  );


  or
  g1655
  (
    n1681,
    n1318,
    n1023,
    n1255,
    n1179
  );


  and
  g1656
  (
    n1670,
    n1212,
    n1342,
    n1099,
    n1334
  );


  or
  g1657
  (
    n1667,
    n1341,
    n1261,
    n1038,
    n1090
  );


  xor
  g1658
  (
    n1625,
    n1276,
    n1322,
    n1132,
    n1313
  );


  xor
  g1659
  (
    n1684,
    n1229,
    n1370,
    n1120,
    n1066
  );


  nand
  g1660
  (
    n1693,
    n1166,
    n1344,
    n1312,
    n1290
  );


  buf
  g1661
  (
    n1713,
    n355
  );


  buf
  g1662
  (
    n1716,
    n1605
  );


  not
  g1663
  (
    n1695,
    n365
  );


  not
  g1664
  (
    n1708,
    n1609
  );


  not
  g1665
  (
    n1724,
    n992
  );


  not
  g1666
  (
    n1717,
    n358
  );


  nor
  g1667
  (
    n1714,
    n354,
    n360
  );


  nand
  g1668
  (
    n1718,
    n990,
    n1610,
    n353,
    n362
  );


  and
  g1669
  (
    n1702,
    n1626,
    n362,
    n1630,
    n358
  );


  xnor
  g1670
  (
    n1698,
    n360,
    n354,
    n364,
    n1614
  );


  nand
  g1671
  (
    n1699,
    n1604,
    n1601,
    n1625,
    n357
  );


  xnor
  g1672
  (
    n1720,
    n364,
    n991,
    n1631,
    n1629
  );


  or
  g1673
  (
    n1709,
    n356,
    n365,
    n355,
    n360
  );


  or
  g1674
  (
    n1700,
    n358,
    n992,
    n991,
    n357
  );


  or
  g1675
  (
    n1711,
    n363,
    n1627,
    n1615,
    n1603
  );


  xor
  g1676
  (
    n1703,
    n1600,
    n1620,
    n357,
    n1622
  );


  or
  g1677
  (
    n1694,
    n356,
    n366,
    n1598,
    n1606
  );


  or
  g1678
  (
    n1715,
    n362,
    n991,
    n1616,
    n1617
  );


  or
  g1679
  (
    n1701,
    n361,
    n1602,
    n357,
    n1612
  );


  or
  g1680
  (
    n1722,
    n1632,
    n991,
    n365,
    n1599
  );


  nand
  g1681
  (
    n1706,
    n364,
    n1618,
    n361,
    n355
  );


  or
  g1682
  (
    n1723,
    n366,
    n1621,
    n358,
    n1619
  );


  nor
  g1683
  (
    n1705,
    n364,
    n990,
    n361,
    n1607
  );


  xor
  g1684
  (
    n1697,
    n1623,
    n363,
    n990,
    n356
  );


  nand
  g1685
  (
    n1719,
    n359,
    n1628,
    n354,
    n366
  );


  xnor
  g1686
  (
    n1696,
    n1613,
    n367,
    n989,
    n366
  );


  or
  g1687
  (
    n1707,
    n355,
    n1634,
    n363,
    n362
  );


  xnor
  g1688
  (
    n1721,
    n1608,
    n363,
    n359
  );


  nand
  g1689
  (
    n1712,
    n361,
    n360,
    n1633,
    n365
  );


  nor
  g1690
  (
    n1704,
    n990,
    n1624,
    n359,
    n367
  );


  nor
  g1691
  (
    n1710,
    n354,
    n1611,
    n356,
    n1635
  );


  and
  g1692
  (
    n1733,
    n1400,
    n1703,
    n1420,
    n1417
  );


  nand
  g1693
  (
    n1734,
    n1394,
    n1416,
    n1396,
    n1701
  );


  xor
  g1694
  (
    n1730,
    n1415,
    n1412,
    n1408,
    n1699
  );


  xnor
  g1695
  (
    n1727,
    n1398,
    n1402,
    n1696,
    n1407
  );


  and
  g1696
  (
    n1731,
    n1418,
    n1700,
    n1419,
    n1697
  );


  xnor
  g1697
  (
    n1726,
    n1405,
    n1393,
    n1414,
    n1403
  );


  and
  g1698
  (
    n1725,
    n1421,
    n1409,
    n1410,
    n1399
  );


  xnor
  g1699
  (
    n1729,
    n1702,
    n1406,
    n1413,
    n1698
  );


  nand
  g1700
  (
    n1732,
    n1694,
    n1422,
    n1395,
    n1397
  );


  xnor
  g1701
  (
    n1728,
    n1411,
    n1695,
    n1401,
    n1404
  );


  nor
  g1702
  (
    n1744,
    n1445,
    n1446,
    n1729,
    n1433
  );


  nand
  g1703
  (
    KeyWire_0_14,
    n1450,
    n1429,
    n1434,
    n1734
  );


  nand
  g1704
  (
    n1735,
    n1727,
    n1423,
    n1430,
    n1442
  );


  or
  g1705
  (
    n1739,
    n1425,
    n1443,
    n1437,
    n1452
  );


  xor
  g1706
  (
    n1745,
    n1432,
    n1441,
    n1436,
    n1428
  );


  nand
  g1707
  (
    n1738,
    n1426,
    n1455,
    n1732,
    n1424
  );


  nand
  g1708
  (
    n1741,
    n1725,
    n1439,
    n1447,
    n1449
  );


  and
  g1709
  (
    n1743,
    n1427,
    n1451,
    n1448,
    n1444
  );


  or
  g1710
  (
    n1742,
    n1728,
    n1440,
    n1431,
    n1731
  );


  nor
  g1711
  (
    n1736,
    n1730,
    n1435,
    n1454,
    n1453
  );


  or
  g1712
  (
    n1737,
    n1734,
    n1726,
    n1438,
    n1733
  );


  nor
  g1713
  (
    n1769,
    n1513,
    n1459,
    n1509,
    n1489
  );


  and
  g1714
  (
    n1774,
    n1490,
    n1542,
    n1494,
    n1739
  );


  xnor
  g1715
  (
    n1758,
    n1506,
    n1492,
    n1499,
    n1735
  );


  nor
  g1716
  (
    n1756,
    n1523,
    n1739,
    n1541,
    n1529
  );


  xnor
  g1717
  (
    n1755,
    n1475,
    n1738,
    n1458,
    n1535
  );


  nor
  g1718
  (
    n1747,
    n1735,
    n1739,
    n1482,
    n1738
  );


  nand
  g1719
  (
    n1751,
    n1740,
    n1486,
    n1484,
    n1736
  );


  nand
  g1720
  (
    n1767,
    n1740,
    n1518,
    n1464,
    n1461
  );


  nor
  g1721
  (
    n1754,
    n1504,
    n1470,
    n1468,
    n1471
  );


  or
  g1722
  (
    n1760,
    n1507,
    n1738,
    n1742,
    n1519
  );


  and
  g1723
  (
    n1763,
    n1525,
    n1480,
    n1737,
    n1500
  );


  nor
  g1724
  (
    n1750,
    n1527,
    n1530,
    n1536,
    n1505
  );


  or
  g1725
  (
    n1761,
    n1545,
    n1456,
    n1520,
    n1462
  );


  xor
  g1726
  (
    n1772,
    n1466,
    n1742,
    n1502,
    n1741
  );


  nor
  g1727
  (
    n1775,
    n1478,
    n1521,
    n1531,
    n1740
  );


  or
  g1728
  (
    n1749,
    n1543,
    n1539,
    n1497,
    n1479
  );


  xnor
  g1729
  (
    n1765,
    n1741,
    n1528,
    n1508,
    n1544
  );


  nand
  g1730
  (
    n1759,
    n1515,
    n1736,
    n1512,
    n1511
  );


  nand
  g1731
  (
    n1773,
    n1460,
    n1737,
    n1501,
    n1487
  );


  or
  g1732
  (
    n1766,
    n1739,
    n1491,
    n1457,
    n1522
  );


  xnor
  g1733
  (
    n1757,
    n1741,
    n1472,
    n1534,
    n1496
  );


  xnor
  g1734
  (
    n1764,
    n1736,
    n1465,
    n1538,
    n1540
  );


  and
  g1735
  (
    n1746,
    n1735,
    n1467,
    n1481,
    n1510
  );


  xor
  g1736
  (
    n1762,
    n1473,
    n1735,
    n1474,
    n1514
  );


  and
  g1737
  (
    n1753,
    n1463,
    n1737,
    n1740,
    n1526
  );


  xor
  g1738
  (
    n1771,
    n1483,
    n1485,
    n1737,
    n1537
  );


  xnor
  g1739
  (
    n1770,
    n1524,
    n1533,
    n1736,
    n1738
  );


  nand
  g1740
  (
    n1768,
    n1503,
    n1477,
    n1476,
    n1495
  );


  or
  g1741
  (
    n1752,
    n1516,
    n1517,
    n1741,
    n1498
  );


  or
  g1742
  (
    n1748,
    n1493,
    n1469,
    n1488,
    n1532
  );


  buf
  g1743
  (
    n1804,
    n1759
  );


  buf
  g1744
  (
    n1777,
    n1751
  );


  not
  g1745
  (
    n1793,
    n1747
  );


  buf
  g1746
  (
    n1813,
    n1747
  );


  not
  g1747
  (
    n1799,
    n1757
  );


  buf
  g1748
  (
    n1789,
    n1749
  );


  buf
  g1749
  (
    n1781,
    n1750
  );


  buf
  g1750
  (
    n1803,
    n1748
  );


  buf
  g1751
  (
    n1800,
    n1756
  );


  buf
  g1752
  (
    n1787,
    n1746
  );


  buf
  g1753
  (
    n1794,
    n1755
  );


  not
  g1754
  (
    n1779,
    n1758
  );


  not
  g1755
  (
    n1807,
    n1749
  );


  not
  g1756
  (
    n1812,
    n1749
  );


  buf
  g1757
  (
    n1814,
    n1746
  );


  buf
  g1758
  (
    n1791,
    n1752
  );


  buf
  g1759
  (
    n1784,
    n1757
  );


  not
  g1760
  (
    n1801,
    n1753
  );


  not
  g1761
  (
    n1776,
    n1757
  );


  not
  g1762
  (
    n1783,
    n1754
  );


  buf
  g1763
  (
    n1802,
    n1755
  );


  not
  g1764
  (
    n1797,
    n1753
  );


  not
  g1765
  (
    n1796,
    n1751
  );


  not
  g1766
  (
    n1810,
    n1751
  );


  not
  g1767
  (
    n1786,
    n1752
  );


  not
  g1768
  (
    n1792,
    n1754
  );


  not
  g1769
  (
    n1798,
    n1759
  );


  buf
  g1770
  (
    n1782,
    n1748
  );


  not
  g1771
  (
    n1811,
    n1750
  );


  not
  g1772
  (
    n1790,
    n1756
  );


  buf
  g1773
  (
    n1788,
    n1747
  );


  buf
  g1774
  (
    n1806,
    n1752
  );


  xor
  g1775
  (
    n1809,
    n1755,
    n1752,
    n1746,
    n1749
  );


  xnor
  g1776
  (
    n1780,
    n1758,
    n1754,
    n1755,
    n1636
  );


  nor
  g1777
  (
    n1795,
    n1751,
    n1754,
    n1756,
    n1758
  );


  and
  g1778
  (
    n1778,
    n1760,
    n1638,
    n1753,
    n1637
  );


  nor
  g1779
  (
    n1808,
    n1750,
    n1759,
    n1753
  );


  nor
  g1780
  (
    n1805,
    n1756,
    n1746,
    n1750,
    n1748
  );


  and
  g1781
  (
    n1785,
    n1757,
    n1758,
    n1747,
    n1748
  );


  and
  g1782
  (
    n1835,
    n994,
    n120,
    n1790,
    n1762
  );


  xor
  g1783
  (
    n1836,
    n1654,
    n1720,
    n1794,
    n1786
  );


  nor
  g1784
  (
    n1820,
    n1717,
    n1783,
    n1554,
    n1558
  );


  or
  g1785
  (
    n1825,
    n1766,
    n1788,
    n1811,
    n1557
  );


  xor
  g1786
  (
    n1839,
    n1791,
    n1646,
    n1807,
    n994
  );


  nand
  g1787
  (
    n1848,
    n1805,
    n55,
    n1799,
    n1707
  );


  xor
  g1788
  (
    n1837,
    n1801,
    n1766,
    n1553,
    n1806
  );


  nand
  g1789
  (
    n1845,
    n1706,
    n1762,
    n1724,
    n1645
  );


  xor
  g1790
  (
    n1831,
    n1710,
    n1813,
    n55,
    n993
  );


  or
  g1791
  (
    n1830,
    n1556,
    n1760,
    n1765,
    n1642
  );


  and
  g1792
  (
    n1822,
    n1718,
    n1715,
    n1640,
    n55
  );


  xnor
  g1793
  (
    n1826,
    n1559,
    n1793,
    n1812,
    n1764
  );


  xor
  g1794
  (
    n1829,
    n1651,
    n1803,
    n1764,
    n1808
  );


  nand
  g1795
  (
    n1843,
    n8,
    n1653,
    n1779,
    n1778
  );


  or
  g1796
  (
    n1850,
    n1644,
    n1814,
    n121,
    n1762
  );


  xor
  g1797
  (
    n1842,
    n121,
    n1760,
    n1782,
    n1797
  );


  xor
  g1798
  (
    n1818,
    n1792,
    n7,
    n1789,
    n994
  );


  nor
  g1799
  (
    n1816,
    n9,
    n120,
    n1764,
    n1709
  );


  xor
  g1800
  (
    n1851,
    n993,
    n1711,
    n1724,
    n9
  );


  nand
  g1801
  (
    n1821,
    n6,
    n992,
    n995,
    n1722
  );


  and
  g1802
  (
    n1827,
    n1649,
    n1763,
    n1765,
    n1814
  );


  nand
  g1803
  (
    n1815,
    n1714,
    n992,
    n1721,
    n1761
  );


  nand
  g1804
  (
    n1834,
    n1704,
    n1648,
    n1712,
    n1776
  );


  xor
  g1805
  (
    n1854,
    n1796,
    n1723,
    n1546,
    n1781
  );


  nor
  g1806
  (
    n1846,
    n119,
    n120,
    n8,
    n1763
  );


  nor
  g1807
  (
    n1853,
    n10,
    n1787,
    n1547,
    n1652
  );


  xnor
  g1808
  (
    n1832,
    n1552,
    n9,
    n1784,
    n1762
  );


  xor
  g1809
  (
    n1841,
    n1764,
    n1802,
    n1647,
    n1763
  );


  nor
  g1810
  (
    n1844,
    n1548,
    n994,
    n1761,
    n995
  );


  or
  g1811
  (
    n1847,
    n7,
    n9,
    n121,
    n1765
  );


  or
  g1812
  (
    n1852,
    n1551,
    n1760,
    n1780,
    n1777
  );


  nor
  g1813
  (
    n1833,
    n1708,
    n7,
    n1639,
    n8
  );


  nor
  g1814
  (
    n1838,
    n1766,
    n10,
    n1763,
    n993
  );


  or
  g1815
  (
    n1824,
    n1810,
    n1785,
    n7,
    n1809
  );


  or
  g1816
  (
    n1819,
    n1555,
    n1804,
    n1761,
    n1550
  );


  or
  g1817
  (
    n1823,
    n1765,
    n1705,
    n1716,
    n8
  );


  nor
  g1818
  (
    n1849,
    n1761,
    n1549,
    n1650,
    n1798
  );


  nor
  g1819
  (
    n1840,
    n1795,
    n1643,
    n1560,
    n995
  );


  nor
  g1820
  (
    n1828,
    n119,
    n993,
    n1641,
    n120
  );


  or
  g1821
  (
    n1817,
    n1719,
    n1713,
    n1800,
    n1561
  );


  not
  g1822
  (
    n1876,
    n1844
  );


  not
  g1823
  (
    n1868,
    n1829
  );


  not
  g1824
  (
    n1874,
    n1838
  );


  buf
  g1825
  (
    n1869,
    n1833
  );


  buf
  g1826
  (
    n1884,
    n1815
  );


  buf
  g1827
  (
    n1860,
    n1840
  );


  not
  g1828
  (
    n1864,
    n1841
  );


  buf
  g1829
  (
    n1855,
    n1834
  );


  buf
  g1830
  (
    n1882,
    n1842
  );


  buf
  g1831
  (
    n1877,
    n1842
  );


  buf
  g1832
  (
    n1859,
    n1830
  );


  buf
  g1833
  (
    n1865,
    n1837
  );


  not
  g1834
  (
    n1871,
    n1845
  );


  buf
  g1835
  (
    n1861,
    n1827
  );


  buf
  g1836
  (
    n1867,
    n1819
  );


  buf
  g1837
  (
    n1872,
    n1826
  );


  not
  g1838
  (
    n1883,
    n1822
  );


  buf
  g1839
  (
    n1873,
    n1821
  );


  not
  g1840
  (
    n1863,
    n1818
  );


  not
  g1841
  (
    n1858,
    n1843
  );


  nand
  g1842
  (
    n1875,
    n1843,
    n1837,
    n1846
  );


  nand
  g1843
  (
    n1881,
    n1838,
    n1836,
    n1824
  );


  or
  g1844
  (
    n1857,
    n1838,
    n1844,
    n1828
  );


  or
  g1845
  (
    n1878,
    n1825,
    n1817,
    n1844
  );


  xor
  g1846
  (
    n1862,
    n1831,
    n1842,
    n1843
  );


  nand
  g1847
  (
    n1856,
    n1835,
    n1836,
    n1832
  );


  xor
  g1848
  (
    n1866,
    n1840,
    n1841,
    n1845
  );


  or
  g1849
  (
    n1880,
    n1841,
    n1845,
    n1823
  );


  xnor
  g1850
  (
    n1879,
    n1820,
    n1836,
    n1837
  );


  or
  g1851
  (
    n1870,
    n1839,
    n1816,
    n1846
  );


  nor
  g1852
  (
    n1885,
    n1846,
    n1840,
    n1839
  );


  and
  g1853
  (
    n1904,
    n1875,
    n1856,
    n1878,
    n15
  );


  and
  g1854
  (
    n1902,
    n24,
    n32,
    n26,
    n10
  );


  and
  g1855
  (
    n1890,
    n1877,
    n31,
    n32,
    n26
  );


  or
  g1856
  (
    n1899,
    n1860,
    n30,
    n1883,
    n17
  );


  xor
  g1857
  (
    n1907,
    n20,
    n1864,
    n29,
    n13
  );


  nand
  g1858
  (
    n1887,
    n27,
    n14,
    n22,
    n1881
  );


  xor
  g1859
  (
    n1908,
    n28,
    n16,
    n20,
    n1855
  );


  xnor
  g1860
  (
    n1906,
    n30,
    n32,
    n19,
    n23
  );


  xnor
  g1861
  (
    n1911,
    n16,
    n31,
    n19,
    n12
  );


  or
  g1862
  (
    n1896,
    n13,
    n11,
    n25,
    n19
  );


  nand
  g1863
  (
    n1912,
    n1874,
    n18,
    n20,
    n29
  );


  and
  g1864
  (
    n1913,
    n13,
    n21,
    n24,
    n1870
  );


  nand
  g1865
  (
    n1903,
    n1882,
    n17,
    n1866
  );


  nand
  g1866
  (
    n1898,
    n16,
    n30,
    n29,
    n1859
  );


  xnor
  g1867
  (
    n1909,
    n15,
    n29,
    n27,
    n22
  );


  and
  g1868
  (
    n1893,
    n1868,
    n28,
    n1861,
    n18
  );


  xor
  g1869
  (
    n1888,
    n10,
    n1869,
    n26,
    n25
  );


  and
  g1870
  (
    n1901,
    n32,
    n1876,
    n13,
    n1880
  );


  xor
  g1871
  (
    n1891,
    n28,
    n14,
    n12,
    n23
  );


  xor
  g1872
  (
    n1895,
    n11,
    n18,
    n24,
    n15
  );


  xor
  g1873
  (
    n1886,
    n25,
    n31,
    n1872,
    n24
  );


  nor
  g1874
  (
    n1897,
    n1862,
    n28,
    n31,
    n12
  );


  nor
  g1875
  (
    n1889,
    n17,
    n1863,
    n21,
    n1865
  );


  or
  g1876
  (
    n1894,
    n1858,
    n15,
    n12,
    n25
  );


  xnor
  g1877
  (
    n1900,
    n23,
    n22,
    n11
  );


  xor
  g1878
  (
    n1910,
    n1879,
    n26,
    n11,
    n18
  );


  nor
  g1879
  (
    n1905,
    n1867,
    n1857,
    n14,
    n1871
  );


  xnor
  g1880
  (
    n1892,
    n20,
    n27,
    n19,
    n30
  );


  nand
  g1881
  (
    n1915,
    n1884,
    n23,
    n27,
    n21
  );


  xnor
  g1882
  (
    n1914,
    n16,
    n21,
    n1873,
    n14
  );


  buf
  g1883
  (
    n1916,
    n1886
  );


  not
  g1884
  (
    n1917,
    n1887
  );


  not
  g1885
  (
    n1921,
    n1917
  );


  not
  g1886
  (
    n1923,
    n1916
  );


  buf
  g1887
  (
    n1922,
    n1916
  );


  buf
  g1888
  (
    n1918,
    n1916
  );


  not
  g1889
  (
    n1920,
    n1916
  );


  not
  g1890
  (
    n1919,
    n1917
  );


  nand
  g1891
  (
    n1925,
    n1923,
    n1848,
    n1921
  );


  nor
  g1892
  (
    n1924,
    n1847,
    n1923,
    n1919
  );


  xor
  g1893
  (
    n1927,
    n1848,
    n1923,
    n1920,
    n1847
  );


  and
  g1894
  (
    n1926,
    n1849,
    n1849,
    n1922,
    n1847
  );


  nor
  g1895
  (
    n1928,
    n1885,
    n1888,
    n1889,
    n1927
  );


  xnor
  g1896
  (
    n1931,
    n1928,
    n190
  );


  xor
  g1897
  (
    n1932,
    n1892,
    n191,
    n190
  );


  xor
  g1898
  (
    n1929,
    n1891,
    n1928,
    n191
  );


  nand
  g1899
  (
    n1930,
    n192,
    n1890,
    n1928,
    n190
  );


  not
  g1900
  (
    n1933,
    n1931
  );


  not
  g1901
  (
    n1936,
    n1930
  );


  buf
  g1902
  (
    n1938,
    n1931
  );


  not
  g1903
  (
    n1939,
    n367
  );


  buf
  g1904
  (
    n1934,
    n1931
  );


  buf
  g1905
  (
    n1935,
    n1930
  );


  not
  g1906
  (
    n1940,
    n1930
  );


  not
  g1907
  (
    n1941,
    n1931
  );


  xnor
  g1908
  (
    n1937,
    n1930,
    n1929
  );


  or
  g1909
  (
    n1943,
    n1934,
    n1006,
    n1002
  );


  xnor
  g1910
  (
    n1947,
    n1005,
    n1002,
    n1936,
    n999
  );


  nand
  g1911
  (
    n1948,
    n996,
    n1936,
    n998,
    n1000
  );


  or
  g1912
  (
    n1950,
    n1001,
    n1005,
    n1003,
    n1933
  );


  nand
  g1913
  (
    n1942,
    n1933,
    n1934,
    n999,
    n1007
  );


  xor
  g1914
  (
    n1957,
    n1004,
    n997,
    n1935
  );


  xor
  g1915
  (
    n1952,
    n1005,
    n998,
    n1001,
    n1936
  );


  nor
  g1916
  (
    n1956,
    n1934,
    n997,
    n1002
  );


  xor
  g1917
  (
    n1944,
    n996,
    n1933,
    n1006,
    n1935
  );


  or
  g1918
  (
    n1946,
    n1936,
    n999,
    n1007,
    n1933
  );


  or
  g1919
  (
    n1949,
    n1003,
    n1004,
    n998,
    n996
  );


  nor
  g1920
  (
    n1955,
    n1003,
    n1002,
    n996,
    n999
  );


  and
  g1921
  (
    n1953,
    n1004,
    n1004,
    n1000,
    n1935
  );


  or
  g1922
  (
    n1951,
    n1007,
    n998,
    n1934,
    n1001
  );


  nand
  g1923
  (
    n1945,
    n1006,
    n995,
    n1003,
    n1001
  );


  nand
  g1924
  (
    n1954,
    n1935,
    n1000,
    n1005
  );


  xor
  g1925
  (
    n1965,
    n1582,
    n1566,
    n1578,
    n1565
  );


  xor
  g1926
  (
    n1962,
    n1564,
    n1953,
    n1571,
    n1585
  );


  xnor
  g1927
  (
    n1958,
    n1572,
    n1951,
    n1563,
    n1584
  );


  nand
  g1928
  (
    n1964,
    n1570,
    n1568,
    n1583,
    n1581
  );


  and
  g1929
  (
    n1960,
    n1567,
    n1562,
    n1950,
    n1569
  );


  or
  g1930
  (
    n1963,
    n1954,
    n1576,
    n1956,
    n1573
  );


  nand
  g1931
  (
    n1961,
    n1579,
    n1952,
    n1575,
    n1957
  );


  xor
  g1932
  (
    n1959,
    n1955,
    n1577,
    n1574,
    n1580
  );


  xnor
  g1933
  (
    n1970,
    n1961,
    n1676,
    n1660,
    n1964
  );


  or
  g1934
  (
    n1971,
    n1962,
    n1963,
    n1678,
    n1965
  );


  and
  g1935
  (
    n1973,
    n1670,
    n1665,
    n1664,
    n1959
  );


  or
  g1936
  (
    n1974,
    n1674,
    n1679,
    n1666,
    n1657
  );


  or
  g1937
  (
    n1968,
    n1680,
    n1669,
    n1681,
    n1668
  );


  xor
  g1938
  (
    n1972,
    n1655,
    n1659,
    n1661,
    n1677
  );


  and
  g1939
  (
    n1966,
    n1675,
    n1960,
    n1672,
    n1662
  );


  xor
  g1940
  (
    n1967,
    n1965,
    n1673,
    n1658,
    n1663
  );


  xnor
  g1941
  (
    n1969,
    n1656,
    n1958,
    n1667,
    n1671
  );


  and
  g1942
  (
    n1978,
    n1590,
    n1972,
    n1932,
    n1591
  );


  nor
  g1943
  (
    n1975,
    n1974,
    n1971,
    n1682,
    n1932
  );


  and
  g1944
  (
    n1976,
    n1586,
    n1973,
    n1932
  );


  nand
  g1945
  (
    n1977,
    n1587,
    n1592,
    n1589,
    n1588
  );


  xor
  g1946
  (
    n1980,
    n1903,
    n1975,
    n1938
  );


  xor
  g1947
  (
    n1979,
    n1905,
    n1937,
    n1975,
    n1912
  );


  xor
  g1948
  (
    n1993,
    n1914,
    n1939,
    n1977
  );


  and
  g1949
  (
    n1984,
    n1902,
    n1897,
    n1894,
    n1898
  );


  nor
  g1950
  (
    n1988,
    n1978,
    n1937,
    n1685,
    n1904
  );


  and
  g1951
  (
    n1985,
    n1938,
    n1913,
    n1977,
    n1976
  );


  xor
  g1952
  (
    n1982,
    n1593,
    n1901,
    n1940,
    n1976
  );


  xnor
  g1953
  (
    n1983,
    n1915,
    n1907,
    n1977,
    n1895
  );


  xor
  g1954
  (
    n1991,
    n1937,
    n1976,
    n1978,
    n1893
  );


  nor
  g1955
  (
    n1994,
    n1899,
    n1940,
    n1900,
    n1977
  );


  or
  g1956
  (
    n1986,
    n1896,
    n1939,
    n1683,
    n1911
  );


  xor
  g1957
  (
    n1990,
    n1975,
    n1906,
    n1940,
    n1686
  );


  or
  g1958
  (
    n1992,
    n1909,
    n1978,
    n1976,
    n1940
  );


  or
  g1959
  (
    n1981,
    n1941,
    n1939,
    n1937,
    n1938
  );


  or
  g1960
  (
    n1989,
    n1941,
    n1975,
    n1908,
    n1684
  );


  nand
  g1961
  (
    n1987,
    n1941,
    n1941,
    n1978,
    n1910
  );


  nand
  g1962
  (
    n2016,
    n1008,
    n1993,
    n1689
  );


  and
  g1963
  (
    n1995,
    n1849,
    n1854,
    n1852,
    n1981
  );


  xor
  g1964
  (
    n2000,
    n368,
    n1851,
    n1743,
    n1595
  );


  or
  g1965
  (
    n2010,
    n369,
    n1992,
    n1852
  );


  xor
  g1966
  (
    n1999,
    n1850,
    n1989,
    n1984,
    n1983
  );


  xor
  g1967
  (
    n2007,
    n1745,
    n1742,
    n368,
    n193
  );


  nand
  g1968
  (
    n2013,
    n1990,
    n1690,
    n1850,
    n1854
  );


  and
  g1969
  (
    n2014,
    n1854,
    n369,
    n1917,
    n1594
  );


  nor
  g1970
  (
    n2008,
    n1853,
    n1007,
    n192,
    n1743
  );


  and
  g1971
  (
    n1998,
    n1744,
    n369,
    n1987,
    n1693
  );


  xnor
  g1972
  (
    n2006,
    n1597,
    n1008,
    n1744,
    n129
  );


  and
  g1973
  (
    n2017,
    n1692,
    n1743,
    n1742,
    n1979
  );


  or
  g1974
  (
    n2005,
    n1917,
    n367,
    n1982,
    n1853
  );


  xnor
  g1975
  (
    n2001,
    n1994,
    n1991,
    n1008,
    n1993
  );


  and
  g1976
  (
    n2012,
    n1853,
    n368,
    n1745,
    n1994
  );


  and
  g1977
  (
    n2009,
    n1986,
    n1743,
    n1851,
    n192
  );


  or
  g1978
  (
    n1997,
    n1850,
    n1994,
    n1691,
    n1688
  );


  or
  g1979
  (
    n2004,
    n369,
    n1854,
    n1008,
    n1744
  );


  xnor
  g1980
  (
    n2002,
    n1993,
    n1853,
    n1687,
    n1745
  );


  xnor
  g1981
  (
    n1996,
    n192,
    n1992,
    n193,
    n1744
  );


  and
  g1982
  (
    n2011,
    n1994,
    n129,
    n1745,
    n1980
  );


  nand
  g1983
  (
    n2015,
    n1985,
    n121,
    n193,
    n1596
  );


  and
  g1984
  (
    n2003,
    n368,
    n193,
    n1988,
    n1851
  );


  nand
  g1985
  (
    n2030,
    n1772,
    n1772,
    n1997,
    n1771
  );


  and
  g1986
  (
    n2029,
    n1773,
    n1774,
    n1769,
    n1768
  );


  xnor
  g1987
  (
    n2019,
    n1767,
    n1770,
    n1769,
    n1766
  );


  xnor
  g1988
  (
    n2032,
    n2009,
    n1773,
    n1767,
    n1768
  );


  nor
  g1989
  (
    n2025,
    n2005,
    n2002,
    n1774,
    n1768
  );


  xnor
  g1990
  (
    n2024,
    n1774,
    n2001,
    n1771,
    n1767
  );


  xnor
  g1991
  (
    n2027,
    n2017,
    n1775,
    n2013,
    n1772
  );


  nand
  g1992
  (
    n2022,
    n1769,
    n1770,
    n2012
  );


  and
  g1993
  (
    n2023,
    n1995,
    n1775,
    n1773,
    n1767
  );


  nor
  g1994
  (
    n2020,
    n2008,
    n2006,
    n1769,
    n1775
  );


  nand
  g1995
  (
    n2021,
    n2016,
    n1996,
    n1998,
    n1772
  );


  nor
  g1996
  (
    n2028,
    n2015,
    n1768,
    n2014,
    n1999
  );


  and
  g1997
  (
    n2018,
    n2003,
    n1774,
    n2007,
    n2010
  );


  nand
  g1998
  (
    n2026,
    n2011,
    n1773,
    n2004,
    n1771
  );


  nor
  g1999
  (
    n2031,
    n1771,
    n1770,
    n1775,
    n2000
  );


  xor
  KeyGate_0_0
  (
    n798,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n837,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n71,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n466,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n276,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n544,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n973,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n493,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n430,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n212,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n520,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n993,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n1054,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n277,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1740,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n192,
    KeyNOTWire_0_15
  );


endmodule


