

module Stat_1456_22_4
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n1152,
  n1149,
  n1145,
  n1160,
  n1157,
  n1167,
  n1150,
  n1148,
  n1155,
  n1159,
  n1163,
  n1143,
  n1158,
  n1161,
  n1146,
  n1151,
  n1190,
  n1180,
  n1178,
  n1191,
  n1486,
  n1485,
  n1483,
  n1484,
  n1479,
  n1481,
  n1480,
  n1482,
  n1478,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;
  output n1152;output n1149;output n1145;output n1160;output n1157;output n1167;output n1150;output n1148;output n1155;output n1159;output n1163;output n1143;output n1158;output n1161;output n1146;output n1151;output n1190;output n1180;output n1178;output n1191;output n1486;output n1485;output n1483;output n1484;output n1479;output n1481;output n1480;output n1482;output n1478;
  wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1144;wire n1147;wire n1153;wire n1154;wire n1156;wire n1162;wire n1164;wire n1165;wire n1166;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1179;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n85,
    n18
  );


  buf
  g1
  (
    n91,
    n4
  );


  not
  g2
  (
    n83,
    n29
  );


  not
  g3
  (
    n47,
    n14
  );


  not
  g4
  (
    n69,
    n30
  );


  buf
  g5
  (
    n123,
    n24
  );


  buf
  g6
  (
    n125,
    n20
  );


  buf
  g7
  (
    n126,
    n20
  );


  not
  g8
  (
    n33,
    n24
  );


  buf
  g9
  (
    n84,
    n15
  );


  not
  g10
  (
    n121,
    n21
  );


  not
  g11
  (
    n53,
    n26
  );


  buf
  g12
  (
    n140,
    n17
  );


  buf
  g13
  (
    n149,
    n9
  );


  not
  g14
  (
    n75,
    n26
  );


  not
  g15
  (
    n136,
    n27
  );


  buf
  g16
  (
    n42,
    n13
  );


  not
  g17
  (
    n72,
    n11
  );


  buf
  g18
  (
    n57,
    n11
  );


  not
  g19
  (
    n120,
    n8
  );


  not
  g20
  (
    n71,
    n2
  );


  buf
  g21
  (
    n137,
    n19
  );


  buf
  g22
  (
    n41,
    n15
  );


  not
  g23
  (
    n32,
    n21
  );


  buf
  g24
  (
    n116,
    n16
  );


  buf
  g25
  (
    n111,
    n18
  );


  buf
  g26
  (
    n133,
    n16
  );


  not
  g27
  (
    n99,
    n29
  );


  buf
  g28
  (
    n94,
    n3
  );


  buf
  g29
  (
    n105,
    n22
  );


  not
  g30
  (
    n117,
    n9
  );


  not
  g31
  (
    n78,
    n22
  );


  not
  g32
  (
    n80,
    n21
  );


  buf
  g33
  (
    n88,
    n3
  );


  buf
  g34
  (
    n58,
    n22
  );


  not
  g35
  (
    n74,
    n6
  );


  not
  g36
  (
    n98,
    n19
  );


  buf
  g37
  (
    n142,
    n26
  );


  buf
  g38
  (
    n51,
    n12
  );


  buf
  g39
  (
    n73,
    n19
  );


  buf
  g40
  (
    n131,
    n3
  );


  not
  g41
  (
    n81,
    n20
  );


  buf
  g42
  (
    n55,
    n2
  );


  buf
  g43
  (
    n77,
    n4
  );


  buf
  g44
  (
    n63,
    n17
  );


  not
  g45
  (
    n79,
    n6
  );


  buf
  g46
  (
    n115,
    n9
  );


  not
  g47
  (
    n122,
    n13
  );


  buf
  g48
  (
    n112,
    n25
  );


  not
  g49
  (
    n31,
    n25
  );


  buf
  g50
  (
    n96,
    n4
  );


  not
  g51
  (
    n86,
    n12
  );


  buf
  g52
  (
    n34,
    n23
  );


  buf
  g53
  (
    n110,
    n3
  );


  not
  g54
  (
    n49,
    n27
  );


  buf
  g55
  (
    n138,
    n18
  );


  not
  g56
  (
    n113,
    n14
  );


  buf
  g57
  (
    n141,
    n8
  );


  not
  g58
  (
    n54,
    n27
  );


  not
  g59
  (
    n124,
    n24
  );


  not
  g60
  (
    n135,
    n23
  );


  not
  g61
  (
    n56,
    n2
  );


  buf
  g62
  (
    n65,
    n1
  );


  buf
  g63
  (
    n37,
    n28
  );


  not
  g64
  (
    n39,
    n14
  );


  not
  g65
  (
    n50,
    n12
  );


  buf
  g66
  (
    n143,
    n1
  );


  buf
  g67
  (
    n119,
    n23
  );


  buf
  g68
  (
    n150,
    n15
  );


  not
  g69
  (
    n107,
    n28
  );


  not
  g70
  (
    n108,
    n21
  );


  not
  g71
  (
    n38,
    n7
  );


  not
  g72
  (
    n36,
    n4
  );


  buf
  g73
  (
    n66,
    n19
  );


  buf
  g74
  (
    n82,
    n23
  );


  buf
  g75
  (
    n114,
    n30
  );


  not
  g76
  (
    n45,
    n11
  );


  not
  g77
  (
    n90,
    n27
  );


  buf
  g78
  (
    n102,
    n18
  );


  not
  g79
  (
    n127,
    n25
  );


  buf
  g80
  (
    n70,
    n7
  );


  buf
  g81
  (
    n106,
    n30
  );


  not
  g82
  (
    n118,
    n17
  );


  not
  g83
  (
    n35,
    n9
  );


  buf
  g84
  (
    n44,
    n1
  );


  buf
  g85
  (
    n147,
    n7
  );


  buf
  g86
  (
    n130,
    n13
  );


  buf
  g87
  (
    n89,
    n28
  );


  buf
  g88
  (
    n103,
    n10
  );


  not
  g89
  (
    n46,
    n5
  );


  not
  g90
  (
    n52,
    n22
  );


  not
  g91
  (
    n97,
    n29
  );


  buf
  g92
  (
    n129,
    n30
  );


  not
  g93
  (
    n109,
    n29
  );


  not
  g94
  (
    n87,
    n6
  );


  buf
  g95
  (
    n132,
    n8
  );


  buf
  g96
  (
    n61,
    n12
  );


  buf
  g97
  (
    n67,
    n13
  );


  buf
  g98
  (
    n146,
    n16
  );


  buf
  g99
  (
    n59,
    n1
  );


  not
  g100
  (
    n48,
    n24
  );


  not
  g101
  (
    n76,
    n2
  );


  buf
  g102
  (
    n95,
    n10
  );


  buf
  g103
  (
    n144,
    n25
  );


  buf
  g104
  (
    n101,
    n10
  );


  buf
  g105
  (
    n93,
    n5
  );


  not
  g106
  (
    n139,
    n14
  );


  not
  g107
  (
    n104,
    n20
  );


  buf
  g108
  (
    n68,
    n16
  );


  buf
  g109
  (
    n60,
    n26
  );


  not
  g110
  (
    n134,
    n5
  );


  buf
  g111
  (
    n64,
    n5
  );


  buf
  g112
  (
    n148,
    n28
  );


  buf
  g113
  (
    n145,
    n11
  );


  not
  g114
  (
    n128,
    n8
  );


  not
  g115
  (
    n40,
    n15
  );


  not
  g116
  (
    n62,
    n6
  );


  buf
  g117
  (
    n43,
    n7
  );


  buf
  g118
  (
    n100,
    n10
  );


  buf
  g119
  (
    n92,
    n17
  );


  buf
  g120
  (
    n194,
    n125
  );


  not
  g121
  (
    n312,
    n149
  );


  buf
  g122
  (
    n599,
    n64
  );


  not
  g123
  (
    n547,
    n126
  );


  not
  g124
  (
    n513,
    n68
  );


  not
  g125
  (
    n487,
    n118
  );


  not
  g126
  (
    n563,
    n100
  );


  buf
  g127
  (
    n390,
    n71
  );


  not
  g128
  (
    n565,
    n95
  );


  buf
  g129
  (
    n450,
    n144
  );


  not
  g130
  (
    n523,
    n104
  );


  not
  g131
  (
    n488,
    n82
  );


  not
  g132
  (
    n460,
    n79
  );


  buf
  g133
  (
    n574,
    n136
  );


  not
  g134
  (
    n417,
    n74
  );


  not
  g135
  (
    n542,
    n41
  );


  buf
  g136
  (
    n242,
    n127
  );


  not
  g137
  (
    n626,
    n132
  );


  buf
  g138
  (
    n454,
    n112
  );


  buf
  g139
  (
    n617,
    n46
  );


  buf
  g140
  (
    n366,
    n140
  );


  buf
  g141
  (
    n174,
    n109
  );


  not
  g142
  (
    n423,
    n72
  );


  not
  g143
  (
    n201,
    n101
  );


  not
  g144
  (
    n316,
    n31
  );


  not
  g145
  (
    n263,
    n132
  );


  buf
  g146
  (
    n573,
    n77
  );


  buf
  g147
  (
    n583,
    n104
  );


  buf
  g148
  (
    n553,
    n115
  );


  buf
  g149
  (
    n234,
    n96
  );


  buf
  g150
  (
    n156,
    n100
  );


  not
  g151
  (
    n256,
    n108
  );


  not
  g152
  (
    n541,
    n37
  );


  buf
  g153
  (
    n385,
    n90
  );


  not
  g154
  (
    n192,
    n122
  );


  buf
  g155
  (
    n216,
    n122
  );


  buf
  g156
  (
    n622,
    n146
  );


  not
  g157
  (
    n623,
    n32
  );


  buf
  g158
  (
    n451,
    n133
  );


  buf
  g159
  (
    n182,
    n69
  );


  not
  g160
  (
    n437,
    n51
  );


  buf
  g161
  (
    n492,
    n77
  );


  not
  g162
  (
    n181,
    n38
  );


  buf
  g163
  (
    n420,
    n58
  );


  not
  g164
  (
    n255,
    n71
  );


  not
  g165
  (
    n502,
    n71
  );


  buf
  g166
  (
    n393,
    n61
  );


  buf
  g167
  (
    n176,
    n128
  );


  not
  g168
  (
    n306,
    n115
  );


  not
  g169
  (
    n435,
    n144
  );


  not
  g170
  (
    n283,
    n42
  );


  not
  g171
  (
    n484,
    n134
  );


  not
  g172
  (
    n318,
    n136
  );


  not
  g173
  (
    n296,
    n129
  );


  not
  g174
  (
    n398,
    n106
  );


  buf
  g175
  (
    n370,
    n69
  );


  not
  g176
  (
    n329,
    n143
  );


  not
  g177
  (
    n239,
    n135
  );


  buf
  g178
  (
    n259,
    n46
  );


  buf
  g179
  (
    n403,
    n63
  );


  not
  g180
  (
    n594,
    n116
  );


  not
  g181
  (
    n151,
    n40
  );


  not
  g182
  (
    n439,
    n64
  );


  buf
  g183
  (
    n200,
    n106
  );


  buf
  g184
  (
    n528,
    n141
  );


  not
  g185
  (
    n543,
    n68
  );


  buf
  g186
  (
    n337,
    n142
  );


  not
  g187
  (
    n466,
    n42
  );


  not
  g188
  (
    n418,
    n147
  );


  not
  g189
  (
    n223,
    n54
  );


  not
  g190
  (
    n533,
    n38
  );


  not
  g191
  (
    n252,
    n108
  );


  buf
  g192
  (
    n374,
    n134
  );


  buf
  g193
  (
    n383,
    n69
  );


  not
  g194
  (
    n470,
    n75
  );


  buf
  g195
  (
    n505,
    n82
  );


  buf
  g196
  (
    n545,
    n127
  );


  not
  g197
  (
    n291,
    n121
  );


  buf
  g198
  (
    n345,
    n65
  );


  not
  g199
  (
    n157,
    n52
  );


  not
  g200
  (
    n554,
    n94
  );


  not
  g201
  (
    n349,
    n83
  );


  not
  g202
  (
    n585,
    n56
  );


  not
  g203
  (
    n445,
    n109
  );


  not
  g204
  (
    n399,
    n121
  );


  not
  g205
  (
    n612,
    n91
  );


  buf
  g206
  (
    n215,
    n145
  );


  not
  g207
  (
    n177,
    n34
  );


  not
  g208
  (
    n355,
    n66
  );


  not
  g209
  (
    n514,
    n120
  );


  buf
  g210
  (
    n520,
    n56
  );


  buf
  g211
  (
    n197,
    n91
  );


  not
  g212
  (
    n534,
    n65
  );


  not
  g213
  (
    n290,
    n93
  );


  not
  g214
  (
    n332,
    n79
  );


  buf
  g215
  (
    n320,
    n39
  );


  buf
  g216
  (
    n361,
    n88
  );


  buf
  g217
  (
    n433,
    n64
  );


  buf
  g218
  (
    n625,
    n103
  );


  not
  g219
  (
    n253,
    n72
  );


  not
  g220
  (
    n524,
    n85
  );


  buf
  g221
  (
    n170,
    n53
  );


  buf
  g222
  (
    n610,
    n118
  );


  not
  g223
  (
    n456,
    n38
  );


  buf
  g224
  (
    n507,
    n60
  );


  not
  g225
  (
    n600,
    n113
  );


  not
  g226
  (
    n568,
    n90
  );


  buf
  g227
  (
    n213,
    n107
  );


  buf
  g228
  (
    n516,
    n45
  );


  not
  g229
  (
    n476,
    n73
  );


  not
  g230
  (
    n331,
    n95
  );


  buf
  g231
  (
    n464,
    n119
  );


  not
  g232
  (
    n493,
    n60
  );


  buf
  g233
  (
    n235,
    n62
  );


  buf
  g234
  (
    n292,
    n117
  );


  not
  g235
  (
    n365,
    n48
  );


  not
  g236
  (
    n159,
    n137
  );


  buf
  g237
  (
    n571,
    n133
  );


  buf
  g238
  (
    n434,
    n95
  );


  not
  g239
  (
    n236,
    n86
  );


  buf
  g240
  (
    n305,
    n34
  );


  buf
  g241
  (
    n472,
    n63
  );


  buf
  g242
  (
    n430,
    n103
  );


  not
  g243
  (
    n188,
    n105
  );


  not
  g244
  (
    n452,
    n80
  );


  not
  g245
  (
    n491,
    n138
  );


  not
  g246
  (
    n604,
    n58
  );


  not
  g247
  (
    n474,
    n32
  );


  not
  g248
  (
    n226,
    n102
  );


  buf
  g249
  (
    n531,
    n137
  );


  buf
  g250
  (
    n480,
    n139
  );


  not
  g251
  (
    n581,
    n47
  );


  buf
  g252
  (
    n247,
    n41
  );


  not
  g253
  (
    n334,
    n98
  );


  not
  g254
  (
    n481,
    n49
  );


  not
  g255
  (
    n429,
    n136
  );


  not
  g256
  (
    n187,
    n78
  );


  buf
  g257
  (
    n501,
    n92
  );


  not
  g258
  (
    n372,
    n116
  );


  buf
  g259
  (
    n229,
    n94
  );


  buf
  g260
  (
    n580,
    n118
  );


  buf
  g261
  (
    n549,
    n48
  );


  not
  g262
  (
    n237,
    n114
  );


  buf
  g263
  (
    n530,
    n63
  );


  not
  g264
  (
    n238,
    n108
  );


  buf
  g265
  (
    n588,
    n42
  );


  buf
  g266
  (
    n288,
    n135
  );


  buf
  g267
  (
    n271,
    n43
  );


  not
  g268
  (
    n478,
    n38
  );


  buf
  g269
  (
    n602,
    n130
  );


  buf
  g270
  (
    n425,
    n149
  );


  buf
  g271
  (
    n473,
    n147
  );


  buf
  g272
  (
    n300,
    n67
  );


  buf
  g273
  (
    n260,
    n150
  );


  not
  g274
  (
    n333,
    n119
  );


  buf
  g275
  (
    n616,
    n79
  );


  not
  g276
  (
    n193,
    n85
  );


  not
  g277
  (
    n232,
    n32
  );


  buf
  g278
  (
    n311,
    n126
  );


  not
  g279
  (
    n392,
    n97
  );


  buf
  g280
  (
    n546,
    n61
  );


  buf
  g281
  (
    n154,
    n124
  );


  buf
  g282
  (
    n397,
    n87
  );


  buf
  g283
  (
    n419,
    n114
  );


  not
  g284
  (
    n576,
    n76
  );


  buf
  g285
  (
    n391,
    n126
  );


  buf
  g286
  (
    n467,
    n147
  );


  buf
  g287
  (
    n338,
    n90
  );


  buf
  g288
  (
    n489,
    n80
  );


  not
  g289
  (
    n225,
    n144
  );


  buf
  g290
  (
    n587,
    n88
  );


  buf
  g291
  (
    n165,
    n68
  );


  not
  g292
  (
    n426,
    n115
  );


  not
  g293
  (
    n497,
    n73
  );


  buf
  g294
  (
    n293,
    n110
  );


  buf
  g295
  (
    n274,
    n61
  );


  buf
  g296
  (
    n586,
    n132
  );


  buf
  g297
  (
    n387,
    n89
  );


  buf
  g298
  (
    n352,
    n68
  );


  not
  g299
  (
    n317,
    n103
  );


  buf
  g300
  (
    n609,
    n96
  );


  buf
  g301
  (
    n195,
    n146
  );


  buf
  g302
  (
    n353,
    n140
  );


  not
  g303
  (
    n526,
    n117
  );


  buf
  g304
  (
    n475,
    n75
  );


  not
  g305
  (
    n308,
    n31
  );


  not
  g306
  (
    n431,
    n141
  );


  buf
  g307
  (
    n540,
    n51
  );


  buf
  g308
  (
    n294,
    n45
  );


  not
  g309
  (
    n369,
    n98
  );


  not
  g310
  (
    n564,
    n139
  );


  not
  g311
  (
    n518,
    n119
  );


  not
  g312
  (
    n506,
    n103
  );


  buf
  g313
  (
    n282,
    n121
  );


  not
  g314
  (
    n438,
    n141
  );


  buf
  g315
  (
    n382,
    n130
  );


  not
  g316
  (
    n619,
    n48
  );


  buf
  g317
  (
    n251,
    n81
  );


  not
  g318
  (
    n499,
    n37
  );


  buf
  g319
  (
    n529,
    n69
  );


  buf
  g320
  (
    n504,
    n97
  );


  not
  g321
  (
    n371,
    n93
  );


  buf
  g322
  (
    n453,
    n90
  );


  buf
  g323
  (
    n327,
    n55
  );


  not
  g324
  (
    n303,
    n65
  );


  not
  g325
  (
    n191,
    n52
  );


  buf
  g326
  (
    n350,
    n42
  );


  buf
  g327
  (
    n198,
    n37
  );


  not
  g328
  (
    n527,
    n112
  );


  not
  g329
  (
    n180,
    n47
  );


  not
  g330
  (
    n572,
    n83
  );


  not
  g331
  (
    n630,
    n120
  );


  buf
  g332
  (
    n249,
    n135
  );


  not
  g333
  (
    n266,
    n119
  );


  buf
  g334
  (
    n627,
    n132
  );


  buf
  g335
  (
    n348,
    n33
  );


  buf
  g336
  (
    n368,
    n31
  );


  not
  g337
  (
    n405,
    n85
  );


  buf
  g338
  (
    n277,
    n44
  );


  buf
  g339
  (
    n449,
    n92
  );


  not
  g340
  (
    n455,
    n150
  );


  buf
  g341
  (
    n440,
    n125
  );


  not
  g342
  (
    n384,
    n97
  );


  not
  g343
  (
    n624,
    n143
  );


  buf
  g344
  (
    n167,
    n111
  );


  not
  g345
  (
    n442,
    n138
  );


  buf
  g346
  (
    n205,
    n87
  );


  not
  g347
  (
    n615,
    n62
  );


  buf
  g348
  (
    n330,
    n147
  );


  not
  g349
  (
    n299,
    n78
  );


  not
  g350
  (
    n284,
    n116
  );


  not
  g351
  (
    n559,
    n79
  );


  not
  g352
  (
    n342,
    n139
  );


  not
  g353
  (
    n519,
    n78
  );


  not
  g354
  (
    n628,
    n130
  );


  not
  g355
  (
    n189,
    n148
  );


  not
  g356
  (
    n539,
    n136
  );


  not
  g357
  (
    n272,
    n124
  );


  not
  g358
  (
    n412,
    n46
  );


  buf
  g359
  (
    n347,
    n143
  );


  buf
  g360
  (
    n544,
    n89
  );


  not
  g361
  (
    n407,
    n61
  );


  buf
  g362
  (
    n560,
    n140
  );


  not
  g363
  (
    n278,
    n126
  );


  not
  g364
  (
    n608,
    n67
  );


  not
  g365
  (
    n386,
    n84
  );


  buf
  g366
  (
    n447,
    n122
  );


  buf
  g367
  (
    n168,
    n131
  );


  buf
  g368
  (
    n289,
    n66
  );


  buf
  g369
  (
    n389,
    n88
  );


  not
  g370
  (
    n269,
    n83
  );


  buf
  g371
  (
    n326,
    n113
  );


  not
  g372
  (
    n307,
    n143
  );


  not
  g373
  (
    n601,
    n105
  );


  not
  g374
  (
    n555,
    n145
  );


  not
  g375
  (
    n315,
    n39
  );


  not
  g376
  (
    n172,
    n47
  );


  buf
  g377
  (
    n413,
    n137
  );


  not
  g378
  (
    n244,
    n48
  );


  not
  g379
  (
    n344,
    n110
  );


  buf
  g380
  (
    n186,
    n72
  );


  buf
  g381
  (
    n185,
    n44
  );


  buf
  g382
  (
    n458,
    n35
  );


  not
  g383
  (
    n522,
    n49
  );


  buf
  g384
  (
    n319,
    n81
  );


  not
  g385
  (
    n336,
    n60
  );


  not
  g386
  (
    n510,
    n142
  );


  not
  g387
  (
    n160,
    n43
  );


  buf
  g388
  (
    n629,
    n36
  );


  not
  g389
  (
    n468,
    n91
  );


  not
  g390
  (
    n376,
    n97
  );


  not
  g391
  (
    n428,
    n88
  );


  not
  g392
  (
    n379,
    n96
  );


  buf
  g393
  (
    n264,
    n142
  );


  not
  g394
  (
    n457,
    n86
  );


  buf
  g395
  (
    n325,
    n144
  );


  not
  g396
  (
    n339,
    n111
  );


  not
  g397
  (
    n508,
    n104
  );


  not
  g398
  (
    n552,
    n87
  );


  buf
  g399
  (
    n551,
    n59
  );


  buf
  g400
  (
    n396,
    n58
  );


  buf
  g401
  (
    n614,
    n114
  );


  not
  g402
  (
    n500,
    n149
  );


  buf
  g403
  (
    n459,
    n123
  );


  buf
  g404
  (
    n550,
    n99
  );


  not
  g405
  (
    n603,
    n118
  );


  not
  g406
  (
    n471,
    n77
  );


  not
  g407
  (
    n377,
    n123
  );


  not
  g408
  (
    n228,
    n112
  );


  buf
  g409
  (
    n286,
    n63
  );


  not
  g410
  (
    n593,
    n123
  );


  buf
  g411
  (
    n224,
    n84
  );


  not
  g412
  (
    n323,
    n53
  );


  not
  g413
  (
    n257,
    n91
  );


  buf
  g414
  (
    n163,
    n124
  );


  not
  g415
  (
    n591,
    n37
  );


  not
  g416
  (
    n482,
    n33
  );


  not
  g417
  (
    n220,
    n81
  );


  buf
  g418
  (
    n394,
    n44
  );


  buf
  g419
  (
    n512,
    n145
  );


  not
  g420
  (
    n485,
    n123
  );


  not
  g421
  (
    n570,
    n100
  );


  not
  g422
  (
    n486,
    n76
  );


  buf
  g423
  (
    n606,
    n39
  );


  not
  g424
  (
    n388,
    n149
  );


  buf
  g425
  (
    n267,
    n67
  );


  not
  g426
  (
    n275,
    n33
  );


  not
  g427
  (
    n321,
    n34
  );


  not
  g428
  (
    n309,
    n54
  );


  not
  g429
  (
    n202,
    n47
  );


  buf
  g430
  (
    n314,
    n82
  );


  not
  g431
  (
    n584,
    n100
  );


  not
  g432
  (
    n184,
    n73
  );


  not
  g433
  (
    n222,
    n80
  );


  not
  g434
  (
    n212,
    n130
  );


  not
  g435
  (
    n246,
    n111
  );


  buf
  g436
  (
    n595,
    n70
  );


  not
  g437
  (
    n313,
    n36
  );


  not
  g438
  (
    n590,
    n138
  );


  buf
  g439
  (
    n178,
    n55
  );


  buf
  g440
  (
    n582,
    n150
  );


  not
  g441
  (
    n569,
    n125
  );


  not
  g442
  (
    n233,
    n92
  );


  not
  g443
  (
    n567,
    n50
  );


  buf
  g444
  (
    n335,
    n117
  );


  buf
  g445
  (
    n532,
    n114
  );


  buf
  g446
  (
    n248,
    n51
  );


  buf
  g447
  (
    n479,
    n141
  );


  buf
  g448
  (
    n561,
    n76
  );


  buf
  g449
  (
    n328,
    n56
  );


  buf
  g450
  (
    n477,
    n109
  );


  not
  g451
  (
    n304,
    n115
  );


  buf
  g452
  (
    n406,
    n148
  );


  buf
  g453
  (
    n175,
    n133
  );


  not
  g454
  (
    n402,
    n36
  );


  buf
  g455
  (
    n621,
    n112
  );


  not
  g456
  (
    n310,
    n57
  );


  not
  g457
  (
    n381,
    n107
  );


  not
  g458
  (
    n556,
    n108
  );


  not
  g459
  (
    n273,
    n117
  );


  buf
  g460
  (
    n268,
    n96
  );


  buf
  g461
  (
    n287,
    n85
  );


  buf
  g462
  (
    n364,
    n84
  );


  not
  g463
  (
    n346,
    n43
  );


  buf
  g464
  (
    n203,
    n59
  );


  buf
  g465
  (
    n432,
    n133
  );


  not
  g466
  (
    n575,
    n107
  );


  not
  g467
  (
    n538,
    n72
  );


  not
  g468
  (
    n153,
    n125
  );


  not
  g469
  (
    n509,
    n120
  );


  not
  g470
  (
    n469,
    n74
  );


  not
  g471
  (
    n483,
    n62
  );


  buf
  g472
  (
    n577,
    n101
  );


  not
  g473
  (
    n265,
    n41
  );


  buf
  g474
  (
    n179,
    n67
  );


  buf
  g475
  (
    n208,
    n146
  );


  buf
  g476
  (
    n162,
    n134
  );


  buf
  g477
  (
    n618,
    n86
  );


  buf
  g478
  (
    n446,
    n50
  );


  not
  g479
  (
    n207,
    n50
  );


  buf
  g480
  (
    n525,
    n138
  );


  buf
  g481
  (
    n262,
    n150
  );


  not
  g482
  (
    n221,
    n129
  );


  not
  g483
  (
    n169,
    n81
  );


  buf
  g484
  (
    n360,
    n131
  );


  not
  g485
  (
    n490,
    n36
  );


  buf
  g486
  (
    n164,
    n105
  );


  not
  g487
  (
    n611,
    n46
  );


  buf
  g488
  (
    n596,
    n52
  );


  not
  g489
  (
    n579,
    n120
  );


  buf
  g490
  (
    n415,
    n102
  );


  buf
  g491
  (
    n199,
    n110
  );


  not
  g492
  (
    n218,
    n93
  );


  buf
  g493
  (
    n562,
    n102
  );


  buf
  g494
  (
    n217,
    n59
  );


  buf
  g495
  (
    n375,
    n32
  );


  not
  g496
  (
    n421,
    n75
  );


  buf
  g497
  (
    n441,
    n116
  );


  not
  g498
  (
    n297,
    n66
  );


  not
  g499
  (
    n322,
    n142
  );


  buf
  g500
  (
    n409,
    n49
  );


  buf
  g501
  (
    n354,
    n148
  );


  not
  g502
  (
    n254,
    n60
  );


  buf
  g503
  (
    n548,
    n129
  );


  buf
  g504
  (
    n359,
    n74
  );


  not
  g505
  (
    n161,
    n75
  );


  buf
  g506
  (
    n589,
    n43
  );


  not
  g507
  (
    n495,
    n57
  );


  not
  g508
  (
    n620,
    n92
  );


  buf
  g509
  (
    n183,
    n52
  );


  not
  g510
  (
    n363,
    n62
  );


  not
  g511
  (
    n152,
    n131
  );


  not
  g512
  (
    n463,
    n148
  );


  buf
  g513
  (
    n400,
    n127
  );


  not
  g514
  (
    n496,
    n86
  );


  not
  g515
  (
    n515,
    n135
  );


  not
  g516
  (
    n408,
    n53
  );


  buf
  g517
  (
    n279,
    n104
  );


  buf
  g518
  (
    n411,
    n95
  );


  not
  g519
  (
    n276,
    n83
  );


  buf
  g520
  (
    n158,
    n131
  );


  not
  g521
  (
    n219,
    n137
  );


  not
  g522
  (
    n285,
    n124
  );


  not
  g523
  (
    n521,
    n44
  );


  not
  g524
  (
    n578,
    n35
  );


  buf
  g525
  (
    n173,
    n84
  );


  not
  g526
  (
    n598,
    n98
  );


  not
  g527
  (
    n416,
    n113
  );


  buf
  g528
  (
    n401,
    n102
  );


  buf
  g529
  (
    n362,
    n34
  );


  buf
  g530
  (
    n231,
    n80
  );


  not
  g531
  (
    n404,
    n146
  );


  buf
  g532
  (
    n414,
    n111
  );


  not
  g533
  (
    n258,
    n70
  );


  buf
  g534
  (
    n607,
    n99
  );


  buf
  g535
  (
    n380,
    n101
  );


  not
  g536
  (
    n324,
    n106
  );


  buf
  g537
  (
    n241,
    n51
  );


  not
  g538
  (
    n613,
    n33
  );


  buf
  g539
  (
    n343,
    n55
  );


  not
  g540
  (
    n295,
    n139
  );


  buf
  g541
  (
    n240,
    n78
  );


  not
  g542
  (
    n461,
    n55
  );


  buf
  g543
  (
    n210,
    n94
  );


  not
  g544
  (
    n357,
    n82
  );


  buf
  g545
  (
    n566,
    n71
  );


  buf
  g546
  (
    n494,
    n99
  );


  buf
  g547
  (
    n281,
    n40
  );


  not
  g548
  (
    n462,
    n59
  );


  buf
  g549
  (
    n503,
    n70
  );


  buf
  g550
  (
    n298,
    n66
  );


  not
  g551
  (
    n261,
    n93
  );


  buf
  g552
  (
    n410,
    n57
  );


  buf
  g553
  (
    n171,
    n64
  );


  buf
  g554
  (
    n302,
    n134
  );


  buf
  g555
  (
    n427,
    n113
  );


  not
  g556
  (
    n245,
    n56
  );


  buf
  g557
  (
    n597,
    n98
  );


  not
  g558
  (
    n230,
    n105
  );


  buf
  g559
  (
    n351,
    n107
  );


  not
  g560
  (
    n448,
    n54
  );


  buf
  g561
  (
    n605,
    n94
  );


  buf
  g562
  (
    n395,
    n53
  );


  buf
  g563
  (
    n517,
    n129
  );


  not
  g564
  (
    n227,
    n35
  );


  not
  g565
  (
    n537,
    n39
  );


  not
  g566
  (
    n211,
    n127
  );


  buf
  g567
  (
    n592,
    n109
  );


  not
  g568
  (
    n204,
    n101
  );


  not
  g569
  (
    n214,
    n49
  );


  not
  g570
  (
    n206,
    n41
  );


  not
  g571
  (
    n422,
    n50
  );


  buf
  g572
  (
    n443,
    n128
  );


  not
  g573
  (
    n301,
    n57
  );


  not
  g574
  (
    n557,
    n65
  );


  buf
  g575
  (
    n558,
    n35
  );


  buf
  g576
  (
    n356,
    n70
  );


  buf
  g577
  (
    n209,
    n54
  );


  buf
  g578
  (
    n373,
    n145
  );


  not
  g579
  (
    n341,
    n76
  );


  buf
  g580
  (
    n358,
    n121
  );


  buf
  g581
  (
    n166,
    n110
  );


  buf
  g582
  (
    n367,
    n128
  );


  not
  g583
  (
    n250,
    n99
  );


  buf
  g584
  (
    n498,
    n31
  );


  not
  g585
  (
    n436,
    n77
  );


  buf
  g586
  (
    n424,
    n58
  );


  not
  g587
  (
    n465,
    n73
  );


  buf
  g588
  (
    n280,
    n45
  );


  not
  g589
  (
    n196,
    n140
  );


  not
  g590
  (
    n511,
    n106
  );


  not
  g591
  (
    n270,
    n89
  );


  not
  g592
  (
    n378,
    n87
  );


  not
  g593
  (
    n340,
    n89
  );


  buf
  g594
  (
    n536,
    n40
  );


  not
  g595
  (
    n155,
    n74
  );


  not
  g596
  (
    n444,
    n128
  );


  buf
  g597
  (
    n535,
    n45
  );


  buf
  g598
  (
    n243,
    n40
  );


  not
  g599
  (
    n190,
    n122
  );


  not
  g600
  (
    n711,
    n429
  );


  buf
  g601
  (
    n659,
    n540
  );


  buf
  g602
  (
    n673,
    n581
  );


  not
  g603
  (
    n725,
    n569
  );


  not
  g604
  (
    n701,
    n565
  );


  buf
  g605
  (
    n690,
    n517
  );


  buf
  g606
  (
    n812,
    n489
  );


  buf
  g607
  (
    n674,
    n530
  );


  buf
  g608
  (
    n683,
    n425
  );


  not
  g609
  (
    n655,
    n403
  );


  not
  g610
  (
    n809,
    n599
  );


  buf
  g611
  (
    n833,
    n428
  );


  buf
  g612
  (
    n756,
    n598
  );


  buf
  g613
  (
    n790,
    n589
  );


  buf
  g614
  (
    n653,
    n577
  );


  buf
  g615
  (
    n767,
    n374
  );


  buf
  g616
  (
    n654,
    n206
  );


  buf
  g617
  (
    n777,
    n584
  );


  not
  g618
  (
    n650,
    n285
  );


  buf
  g619
  (
    n672,
    n407
  );


  not
  g620
  (
    n847,
    n582
  );


  buf
  g621
  (
    n840,
    n344
  );


  buf
  g622
  (
    n752,
    n188
  );


  buf
  g623
  (
    n631,
    n594
  );


  not
  g624
  (
    n783,
    n256
  );


  not
  g625
  (
    n730,
    n616
  );


  buf
  g626
  (
    n676,
    n571
  );


  not
  g627
  (
    n731,
    n388
  );


  buf
  g628
  (
    n667,
    n603
  );


  buf
  g629
  (
    n738,
    n347
  );


  not
  g630
  (
    n838,
    n300
  );


  not
  g631
  (
    n856,
    n595
  );


  not
  g632
  (
    n825,
    n503
  );


  buf
  g633
  (
    n710,
    n611
  );


  not
  g634
  (
    n639,
    n328
  );


  not
  g635
  (
    n721,
    n579
  );


  buf
  g636
  (
    n751,
    n225
  );


  buf
  g637
  (
    n764,
    n524
  );


  buf
  g638
  (
    n824,
    n588
  );


  buf
  g639
  (
    n708,
    n578
  );


  buf
  g640
  (
    n703,
    n368
  );


  not
  g641
  (
    n724,
    n571
  );


  buf
  g642
  (
    n806,
    n596
  );


  buf
  g643
  (
    n677,
    n611
  );


  not
  g644
  (
    n645,
    n358
  );


  not
  g645
  (
    n728,
    n467
  );


  buf
  g646
  (
    n662,
    n313
  );


  not
  g647
  (
    n776,
    n333
  );


  not
  g648
  (
    n827,
    n158
  );


  buf
  g649
  (
    n800,
    n607
  );


  buf
  g650
  (
    n808,
    n377
  );


  not
  g651
  (
    n675,
    n394
  );


  buf
  g652
  (
    n739,
    n601
  );


  not
  g653
  (
    n814,
    n583
  );


  not
  g654
  (
    n831,
    n564
  );


  buf
  g655
  (
    n765,
    n525
  );


  not
  g656
  (
    n671,
    n596
  );


  not
  g657
  (
    n743,
    n537
  );


  not
  g658
  (
    n805,
    n172
  );


  not
  g659
  (
    n795,
    n533
  );


  not
  g660
  (
    n770,
    n568
  );


  not
  g661
  (
    n682,
    n276
  );


  buf
  g662
  (
    n784,
    n608
  );


  not
  g663
  (
    n737,
    n194
  );


  not
  g664
  (
    n759,
    n224
  );


  buf
  g665
  (
    n718,
    n610
  );


  not
  g666
  (
    n702,
    n491
  );


  not
  g667
  (
    n766,
    n557
  );


  buf
  g668
  (
    n664,
    n418
  );


  not
  g669
  (
    n684,
    n519
  );


  buf
  g670
  (
    n757,
    n573
  );


  not
  g671
  (
    n722,
    n463
  );


  not
  g672
  (
    n844,
    n474
  );


  buf
  g673
  (
    n816,
    n461
  );


  not
  g674
  (
    n828,
    n325
  );


  buf
  g675
  (
    n712,
    n528
  );


  not
  g676
  (
    n632,
    n360
  );


  not
  g677
  (
    n758,
    n160
  );


  not
  g678
  (
    n782,
    n550
  );


  buf
  g679
  (
    n697,
    n273
  );


  not
  g680
  (
    n748,
    n547
  );


  buf
  g681
  (
    n747,
    n496
  );


  not
  g682
  (
    n791,
    n342
  );


  not
  g683
  (
    n772,
    n209
  );


  not
  g684
  (
    n678,
    n611
  );


  buf
  g685
  (
    n802,
    n611
  );


  not
  g686
  (
    n850,
    n575
  );


  not
  g687
  (
    n804,
    n471
  );


  buf
  g688
  (
    n637,
    n576
  );


  buf
  g689
  (
    n635,
    n312
  );


  not
  g690
  (
    n796,
    n436
  );


  not
  g691
  (
    n733,
    n364
  );


  nand
  g692
  (
    n723,
    n608,
    n606
  );


  nor
  g693
  (
    n648,
    n258,
    n576
  );


  nor
  g694
  (
    n666,
    n579,
    n161,
    n434,
    n168
  );


  xnor
  g695
  (
    n694,
    n606,
    n290,
    n544,
    n589
  );


  or
  g696
  (
    n842,
    n586,
    n614,
    n581,
    n165
  );


  or
  g697
  (
    n803,
    n598,
    n151,
    n574,
    n326
  );


  xor
  g698
  (
    n686,
    n614,
    n399,
    n171,
    n602
  );


  nor
  g699
  (
    n726,
    n514,
    n581,
    n584,
    n424
  );


  nand
  g700
  (
    n818,
    n350,
    n401,
    n451,
    n597
  );


  nor
  g701
  (
    n636,
    n234,
    n580,
    n462,
    n180
  );


  xnor
  g702
  (
    n736,
    n346,
    n379,
    n588,
    n330
  );


  and
  g703
  (
    n691,
    n204,
    n322,
    n505,
    n438
  );


  or
  g704
  (
    n644,
    n365,
    n526,
    n532,
    n586
  );


  and
  g705
  (
    n741,
    n354,
    n408,
    n602,
    n299
  );


  xnor
  g706
  (
    n778,
    n477,
    n210,
    n417,
    n376
  );


  or
  g707
  (
    n837,
    n187,
    n523,
    n594,
    n269
  );


  or
  g708
  (
    n696,
    n252,
    n192,
    n198,
    n578
  );


  or
  g709
  (
    n661,
    n500,
    n439,
    n534,
    n207
  );


  nor
  g710
  (
    n707,
    n574,
    n405,
    n582,
    n497
  );


  or
  g711
  (
    n641,
    n288,
    n599,
    n179,
    n284
  );


  xor
  g712
  (
    n832,
    n267,
    n321,
    n565,
    n599
  );


  or
  g713
  (
    n642,
    n604,
    n566,
    n185,
    n587
  );


  xor
  g714
  (
    n685,
    n542,
    n308,
    n608,
    n295
  );


  and
  g715
  (
    n769,
    n297,
    n478,
    n591,
    n223
  );


  xnor
  g716
  (
    n815,
    n585,
    n469,
    n603,
    n395
  );


  xnor
  g717
  (
    n775,
    n510,
    n189,
    n375,
    n262
  );


  or
  g718
  (
    n797,
    n522,
    n615,
    n244,
    n466
  );


  nand
  g719
  (
    n735,
    n442,
    n601,
    n255,
    n215
  );


  xnor
  g720
  (
    n760,
    n402,
    n404,
    n603,
    n199
  );


  xnor
  g721
  (
    n660,
    n575,
    n293,
    n304,
    n597
  );


  xor
  g722
  (
    n679,
    n592,
    n574,
    n576,
    n378
  );


  nor
  g723
  (
    n848,
    n334,
    n612,
    n250,
    n575
  );


  nand
  g724
  (
    n633,
    n590,
    n593,
    n162,
    n585
  );


  nor
  g725
  (
    n729,
    n420,
    n373,
    n468,
    n353
  );


  and
  g726
  (
    n755,
    n246,
    n396,
    n298,
    n570
  );


  nor
  g727
  (
    n843,
    n575,
    n421,
    n490,
    n264
  );


  xor
  g728
  (
    n704,
    n578,
    n191,
    n433,
    n613
  );


  and
  g729
  (
    n857,
    n608,
    n459,
    n176,
    n609
  );


  xor
  g730
  (
    n698,
    n564,
    n592,
    n317,
    n566
  );


  nand
  g731
  (
    n792,
    n614,
    n164,
    n260,
    n232
  );


  xor
  g732
  (
    n822,
    n507,
    n535,
    n487,
    n218
  );


  nand
  g733
  (
    n851,
    n338,
    n380,
    n302,
    n600
  );


  nor
  g734
  (
    n788,
    n278,
    n253,
    n190,
    n615
  );


  nor
  g735
  (
    n689,
    n393,
    n612,
    n254,
    n602
  );


  nand
  g736
  (
    n794,
    n183,
    n343,
    n181,
    n348
  );


  or
  g737
  (
    n709,
    n398,
    n577,
    n458,
    n307
  );


  and
  g738
  (
    n719,
    n319,
    n327,
    n597,
    n386
  );


  nor
  g739
  (
    n762,
    n314,
    n247,
    n248,
    n332
  );


  nand
  g740
  (
    n663,
    n239,
    n296,
    n170,
    n242
  );


  or
  g741
  (
    n823,
    n586,
    n320,
    n602,
    n538
  );


  nor
  g742
  (
    n681,
    n283,
    n275,
    n266,
    n559
  );


  xnor
  g743
  (
    n853,
    n587,
    n361,
    n221,
    n583
  );


  xnor
  g744
  (
    n835,
    n549,
    n529,
    n515,
    n201
  );


  and
  g745
  (
    n742,
    n449,
    n460,
    n554,
    n270
  );


  nor
  g746
  (
    n852,
    n511,
    n512,
    n580,
    n592
  );


  xor
  g747
  (
    n658,
    n229,
    n587,
    n567,
    n499
  );


  xnor
  g748
  (
    n830,
    n286,
    n324,
    n289,
    n415
  );


  xnor
  g749
  (
    n716,
    n605,
    n318,
    n222,
    n539
  );


  nand
  g750
  (
    n813,
    n261,
    n167,
    n184,
    n485
  );


  or
  g751
  (
    n705,
    n277,
    n579,
    n600,
    n272
  );


  nand
  g752
  (
    n780,
    n445,
    n588,
    n381,
    n235
  );


  and
  g753
  (
    n798,
    n598,
    n594,
    n603,
    n309
  );


  xnor
  g754
  (
    n829,
    n455,
    n480,
    n166,
    n483
  );


  nand
  g755
  (
    n773,
    n383,
    n454,
    n263,
    n594
  );


  xor
  g756
  (
    n763,
    n169,
    n572,
    n306,
    n589
  );


  xor
  g757
  (
    n670,
    n163,
    n400,
    n280,
    n447
  );


  nand
  g758
  (
    n807,
    n600,
    n614,
    n605,
    n484
  );


  or
  g759
  (
    n669,
    n604,
    n453,
    n612,
    n193
  );


  nor
  g760
  (
    n727,
    n230,
    n504,
    n569,
    n591
  );


  nor
  g761
  (
    n793,
    n574,
    n279,
    n366,
    n563
  );


  xnor
  g762
  (
    n854,
    n352,
    n585,
    n607,
    n593
  );


  and
  g763
  (
    n754,
    n609,
    n212,
    n173,
    n231
  );


  or
  g764
  (
    n799,
    n520,
    n274,
    n493,
    n268
  );


  or
  g765
  (
    n820,
    n432,
    n426,
    n337,
    n604
  );


  or
  g766
  (
    n768,
    n598,
    n572,
    n583,
    n464
  );


  and
  g767
  (
    n692,
    n363,
    n427,
    n152,
    n444
  );


  xnor
  g768
  (
    n634,
    n281,
    n613,
    n456,
    n572
  );


  xnor
  g769
  (
    n753,
    n488,
    n570,
    n572,
    n612
  );


  and
  g770
  (
    n836,
    n349,
    n294,
    n227,
    n174
  );


  xor
  g771
  (
    n810,
    n518,
    n610,
    n582,
    n336
  );


  nand
  g772
  (
    n841,
    n291,
    n605,
    n323,
    n588
  );


  nor
  g773
  (
    n657,
    n331,
    n430,
    n607,
    n546
  );


  nand
  g774
  (
    n855,
    n573,
    n570,
    n521,
    n560
  );


  or
  g775
  (
    n643,
    n531,
    n578,
    n271,
    n335
  );


  nand
  g776
  (
    n845,
    n555,
    n370,
    n516,
    n203
  );


  and
  g777
  (
    n821,
    n482,
    n616,
    n551,
    n583
  );


  or
  g778
  (
    n665,
    n303,
    n384,
    n567,
    n441
  );


  and
  g779
  (
    n668,
    n265,
    n601,
    n566,
    n443
  );


  xor
  g780
  (
    n811,
    n569,
    n566,
    n355,
    n153
  );


  xor
  g781
  (
    n745,
    n568,
    n372,
    n316,
    n177
  );


  nor
  g782
  (
    n706,
    n470,
    n431,
    n205,
    n479
  );


  nor
  g783
  (
    n680,
    n369,
    n553,
    n563,
    n195
  );


  xnor
  g784
  (
    n638,
    n340,
    n481,
    n213,
    n591
  );


  xnor
  g785
  (
    n771,
    n437,
    n413,
    n200,
    n241
  );


  and
  g786
  (
    n720,
    n214,
    n202,
    n564,
    n410
  );


  nand
  g787
  (
    n688,
    n590,
    n576,
    n216,
    n238
  );


  xnor
  g788
  (
    n750,
    n236,
    n584,
    n592,
    n616
  );


  xor
  g789
  (
    n781,
    n411,
    n259,
    n590,
    n541
  );


  nand
  g790
  (
    n819,
    n586,
    n292,
    n389,
    n615
  );


  xnor
  g791
  (
    n789,
    n157,
    n498,
    n552,
    n495
  );


  and
  g792
  (
    n839,
    n604,
    n182,
    n387,
    n513
  );


  and
  g793
  (
    n849,
    n351,
    n208,
    n600,
    n606
  );


  xnor
  g794
  (
    n715,
    n448,
    n567,
    n465,
    n568
  );


  nand
  g795
  (
    n826,
    n607,
    n409,
    n412,
    n573
  );


  nor
  g796
  (
    n732,
    n356,
    n249,
    n509,
    n585
  );


  nand
  g797
  (
    n774,
    n565,
    n186,
    n610,
    n589
  );


  nor
  g798
  (
    n846,
    n579,
    n341,
    n226,
    n301
  );


  xnor
  g799
  (
    n717,
    n345,
    n457,
    n473,
    n220
  );


  xnor
  g800
  (
    n649,
    n217,
    n251,
    n486,
    n587
  );


  xor
  g801
  (
    n785,
    n435,
    n237,
    n536,
    n197
  );


  and
  g802
  (
    n656,
    n414,
    n219,
    n543,
    n423
  );


  nand
  g803
  (
    n695,
    n450,
    n282,
    n371,
    n610
  );


  or
  g804
  (
    n651,
    n367,
    n154,
    n580,
    n595
  );


  xor
  g805
  (
    n746,
    n452,
    n563,
    n556,
    n245
  );


  xnor
  g806
  (
    n713,
    n315,
    n243,
    n545,
    n385
  );


  and
  g807
  (
    n786,
    n502,
    n613,
    n616,
    n582
  );


  xor
  g808
  (
    n779,
    n311,
    n228,
    n595,
    n196
  );


  or
  g809
  (
    n646,
    n590,
    n211,
    n567,
    n175
  );


  xor
  g810
  (
    n817,
    n382,
    n329,
    n584,
    n240
  );


  xnor
  g811
  (
    n714,
    n159,
    n391,
    n606,
    n446
  );


  or
  g812
  (
    n699,
    n416,
    n569,
    n494,
    n476
  );


  nand
  g813
  (
    n734,
    n506,
    n595,
    n571,
    n508
  );


  nor
  g814
  (
    n687,
    n362,
    n605,
    n581,
    n596
  );


  nor
  g815
  (
    n640,
    n178,
    n609,
    n571
  );


  xnor
  g816
  (
    n744,
    n357,
    n422,
    n565,
    n501
  );


  nand
  g817
  (
    n740,
    n564,
    n287,
    n156,
    n233
  );


  xnor
  g818
  (
    n700,
    n472,
    n580,
    n406,
    n390
  );


  nand
  g819
  (
    n787,
    n577,
    n339,
    n527,
    n601
  );


  or
  g820
  (
    n693,
    n155,
    n359,
    n596,
    n597
  );


  nor
  g821
  (
    n647,
    n570,
    n475,
    n492,
    n257
  );


  nand
  g822
  (
    n834,
    n392,
    n615,
    n563,
    n568
  );


  or
  g823
  (
    n761,
    n305,
    n613,
    n440,
    n562
  );


  nand
  g824
  (
    n749,
    n310,
    n419,
    n397,
    n593
  );


  or
  g825
  (
    n652,
    n558,
    n599,
    n593,
    n577
  );


  or
  g826
  (
    n801,
    n548,
    n561,
    n591,
    n573
  );


  buf
  g827
  (
    n917,
    n730
  );


  not
  g828
  (
    n983,
    n682
  );


  buf
  g829
  (
    n947,
    n822
  );


  not
  g830
  (
    n934,
    n805
  );


  buf
  g831
  (
    n1038,
    n850
  );


  buf
  g832
  (
    n1060,
    n842
  );


  not
  g833
  (
    n866,
    n638
  );


  not
  g834
  (
    n1046,
    n845
  );


  buf
  g835
  (
    n982,
    n747
  );


  not
  g836
  (
    n1007,
    n851
  );


  buf
  g837
  (
    n1002,
    n676
  );


  buf
  g838
  (
    n1009,
    n852
  );


  buf
  g839
  (
    n886,
    n748
  );


  not
  g840
  (
    n858,
    n658
  );


  buf
  g841
  (
    n949,
    n820
  );


  buf
  g842
  (
    n930,
    n666
  );


  buf
  g843
  (
    n1040,
    n798
  );


  not
  g844
  (
    n936,
    n818
  );


  buf
  g845
  (
    n990,
    n704
  );


  buf
  g846
  (
    n1013,
    n761
  );


  not
  g847
  (
    n888,
    n819
  );


  buf
  g848
  (
    n887,
    n844
  );


  buf
  g849
  (
    n912,
    n703
  );


  not
  g850
  (
    n1041,
    n722
  );


  not
  g851
  (
    n869,
    n671
  );


  buf
  g852
  (
    n873,
    n802
  );


  buf
  g853
  (
    n879,
    n632
  );


  buf
  g854
  (
    n1044,
    n824
  );


  buf
  g855
  (
    n958,
    n661
  );


  buf
  g856
  (
    n1059,
    n825
  );


  not
  g857
  (
    n968,
    n755
  );


  not
  g858
  (
    n909,
    n795
  );


  not
  g859
  (
    n979,
    n690
  );


  buf
  g860
  (
    n975,
    n815
  );


  not
  g861
  (
    n1000,
    n648
  );


  not
  g862
  (
    n1010,
    n738
  );


  buf
  g863
  (
    n1029,
    n721
  );


  buf
  g864
  (
    n981,
    n830
  );


  not
  g865
  (
    n905,
    n847
  );


  buf
  g866
  (
    n1011,
    n734
  );


  not
  g867
  (
    n1064,
    n712
  );


  buf
  g868
  (
    n1074,
    n735
  );


  not
  g869
  (
    n1052,
    n856
  );


  not
  g870
  (
    n903,
    n760
  );


  not
  g871
  (
    n1061,
    n853
  );


  not
  g872
  (
    n1025,
    n660
  );


  buf
  g873
  (
    n1056,
    n708
  );


  buf
  g874
  (
    n1012,
    n634
  );


  buf
  g875
  (
    n883,
    n695
  );


  not
  g876
  (
    n963,
    n749
  );


  buf
  g877
  (
    n971,
    n736
  );


  not
  g878
  (
    n878,
    n831
  );


  buf
  g879
  (
    n867,
    n793
  );


  not
  g880
  (
    n1039,
    n644
  );


  not
  g881
  (
    n954,
    n724
  );


  not
  g882
  (
    n1032,
    n697
  );


  buf
  g883
  (
    n996,
    n796
  );


  not
  g884
  (
    n948,
    n742
  );


  buf
  g885
  (
    n997,
    n803
  );


  buf
  g886
  (
    n870,
    n836
  );


  buf
  g887
  (
    n1083,
    n709
  );


  buf
  g888
  (
    n980,
    n719
  );


  buf
  g889
  (
    n974,
    n751
  );


  not
  g890
  (
    n1035,
    n698
  );


  not
  g891
  (
    n1062,
    n854
  );


  buf
  g892
  (
    n985,
    n771
  );


  buf
  g893
  (
    n966,
    n725
  );


  buf
  g894
  (
    n942,
    n789
  );


  buf
  g895
  (
    n1045,
    n826
  );


  not
  g896
  (
    n1066,
    n669
  );


  not
  g897
  (
    n976,
    n855
  );


  buf
  g898
  (
    n861,
    n727
  );


  buf
  g899
  (
    n1072,
    n733
  );


  not
  g900
  (
    n1020,
    n776
  );


  not
  g901
  (
    n896,
    n762
  );


  buf
  g902
  (
    n868,
    n678
  );


  not
  g903
  (
    n973,
    n649
  );


  not
  g904
  (
    n892,
    n681
  );


  not
  g905
  (
    n964,
    n821
  );


  buf
  g906
  (
    n956,
    n809
  );


  buf
  g907
  (
    n998,
    n745
  );


  not
  g908
  (
    n961,
    n685
  );


  buf
  g909
  (
    n1075,
    n813
  );


  buf
  g910
  (
    n1003,
    n816
  );


  buf
  g911
  (
    n999,
    n780
  );


  not
  g912
  (
    n984,
    n663
  );


  buf
  g913
  (
    n922,
    n750
  );


  buf
  g914
  (
    n877,
    n715
  );


  not
  g915
  (
    n894,
    n846
  );


  not
  g916
  (
    n863,
    n827
  );


  buf
  g917
  (
    n915,
    n700
  );


  buf
  g918
  (
    n923,
    n645
  );


  not
  g919
  (
    n1008,
    n791
  );


  buf
  g920
  (
    n881,
    n668
  );


  not
  g921
  (
    n913,
    n646
  );


  buf
  g922
  (
    n871,
    n675
  );


  buf
  g923
  (
    n1053,
    n848
  );


  not
  g924
  (
    n926,
    n639
  );


  not
  g925
  (
    n944,
    n804
  );


  buf
  g926
  (
    n957,
    n731
  );


  not
  g927
  (
    n952,
    n792
  );


  buf
  g928
  (
    n972,
    n838
  );


  buf
  g929
  (
    n1005,
    n732
  );


  not
  g930
  (
    n1073,
    n688
  );


  buf
  g931
  (
    n1024,
    n783
  );


  buf
  g932
  (
    n1006,
    n808
  );


  not
  g933
  (
    n938,
    n757
  );


  not
  g934
  (
    n1058,
    n834
  );


  not
  g935
  (
    n1055,
    n806
  );


  not
  g936
  (
    n987,
    n794
  );


  buf
  g937
  (
    n951,
    n758
  );


  not
  g938
  (
    n988,
    n654
  );


  buf
  g939
  (
    n898,
    n728
  );


  not
  g940
  (
    n860,
    n833
  );


  not
  g941
  (
    n885,
    n832
  );


  not
  g942
  (
    n1022,
    n781
  );


  not
  g943
  (
    n910,
    n746
  );


  buf
  g944
  (
    n941,
    n790
  );


  not
  g945
  (
    n1027,
    n829
  );


  buf
  g946
  (
    n906,
    n662
  );


  buf
  g947
  (
    n1068,
    n843
  );


  not
  g948
  (
    n955,
    n674
  );


  buf
  g949
  (
    n1023,
    n782
  );


  not
  g950
  (
    n1065,
    n665
  );


  buf
  g951
  (
    n969,
    n784
  );


  not
  g952
  (
    n932,
    n811
  );


  buf
  g953
  (
    n1026,
    n652
  );


  buf
  g954
  (
    n994,
    n693
  );


  buf
  g955
  (
    n939,
    n786
  );


  buf
  g956
  (
    n1043,
    n759
  );


  not
  g957
  (
    n897,
    n714
  );


  buf
  g958
  (
    n943,
    n655
  );


  not
  g959
  (
    n876,
    n729
  );


  not
  g960
  (
    n1069,
    n707
  );


  buf
  g961
  (
    n1076,
    n810
  );


  not
  g962
  (
    n1019,
    n637
  );


  buf
  g963
  (
    n995,
    n640
  );


  buf
  g964
  (
    n895,
    n679
  );


  not
  g965
  (
    n946,
    n817
  );


  buf
  g966
  (
    n916,
    n683
  );


  not
  g967
  (
    n1081,
    n633
  );


  buf
  g968
  (
    n890,
    n754
  );


  not
  g969
  (
    n978,
    n672
  );


  buf
  g970
  (
    n1057,
    n772
  );


  not
  g971
  (
    n1082,
    n756
  );


  not
  g972
  (
    n924,
    n723
  );


  buf
  g973
  (
    n993,
    n814
  );


  not
  g974
  (
    n1078,
    n774
  );


  buf
  g975
  (
    n1016,
    n694
  );


  not
  g976
  (
    n959,
    n689
  );


  buf
  g977
  (
    n884,
    n686
  );


  not
  g978
  (
    n1036,
    n765
  );


  not
  g979
  (
    n874,
    n785
  );


  not
  g980
  (
    n907,
    n841
  );


  not
  g981
  (
    n1067,
    n764
  );


  buf
  g982
  (
    n962,
    n710
  );


  not
  g983
  (
    n859,
    n677
  );


  not
  g984
  (
    n1054,
    n770
  );


  not
  g985
  (
    n967,
    n769
  );


  not
  g986
  (
    n911,
    n788
  );


  buf
  g987
  (
    n1063,
    n741
  );


  not
  g988
  (
    n1049,
    n777
  );


  buf
  g989
  (
    n960,
    n807
  );


  not
  g990
  (
    n945,
    n839
  );


  not
  g991
  (
    n900,
    n711
  );


  not
  g992
  (
    n901,
    n787
  );


  buf
  g993
  (
    n893,
    n726
  );


  buf
  g994
  (
    n989,
    n837
  );


  buf
  g995
  (
    n872,
    n706
  );


  not
  g996
  (
    n950,
    n647
  );


  buf
  g997
  (
    n1047,
    n642
  );


  buf
  g998
  (
    n921,
    n699
  );


  not
  g999
  (
    n918,
    n739
  );


  buf
  g1000
  (
    n1050,
    n823
  );


  buf
  g1001
  (
    n904,
    n849
  );


  not
  g1002
  (
    n899,
    n656
  );


  not
  g1003
  (
    n935,
    n705
  );


  not
  g1004
  (
    n940,
    n650
  );


  buf
  g1005
  (
    n889,
    n702
  );


  not
  g1006
  (
    n1079,
    n766
  );


  buf
  g1007
  (
    n933,
    n701
  );


  not
  g1008
  (
    n1017,
    n775
  );


  buf
  g1009
  (
    n1030,
    n763
  );


  buf
  g1010
  (
    n1034,
    n744
  );


  not
  g1011
  (
    n908,
    n713
  );


  buf
  g1012
  (
    n929,
    n636
  );


  buf
  g1013
  (
    n1042,
    n653
  );


  buf
  g1014
  (
    n1080,
    n779
  );


  buf
  g1015
  (
    n1004,
    n740
  );


  not
  g1016
  (
    n1037,
    n800
  );


  not
  g1017
  (
    n1071,
    n657
  );


  buf
  g1018
  (
    n977,
    n812
  );


  not
  g1019
  (
    n1018,
    n737
  );


  buf
  g1020
  (
    n991,
    n667
  );


  buf
  g1021
  (
    n875,
    n684
  );


  not
  g1022
  (
    n1031,
    n828
  );


  buf
  g1023
  (
    n1048,
    n720
  );


  not
  g1024
  (
    n1028,
    n797
  );


  buf
  g1025
  (
    n931,
    n631
  );


  not
  g1026
  (
    n925,
    n799
  );


  buf
  g1027
  (
    n914,
    n840
  );


  not
  g1028
  (
    n902,
    n687
  );


  buf
  g1029
  (
    n1021,
    n673
  );


  buf
  g1030
  (
    n965,
    n753
  );


  buf
  g1031
  (
    n891,
    n641
  );


  not
  g1032
  (
    n864,
    n651
  );


  not
  g1033
  (
    n1014,
    n801
  );


  buf
  g1034
  (
    n953,
    n717
  );


  buf
  g1035
  (
    n1077,
    n664
  );


  not
  g1036
  (
    n1001,
    n835
  );


  buf
  g1037
  (
    n882,
    n691
  );


  not
  g1038
  (
    n927,
    n659
  );


  buf
  g1039
  (
    n880,
    n768
  );


  not
  g1040
  (
    n865,
    n696
  );


  not
  g1041
  (
    n1015,
    n752
  );


  buf
  g1042
  (
    n937,
    n767
  );


  buf
  g1043
  (
    n1051,
    n635
  );


  not
  g1044
  (
    n986,
    n716
  );


  buf
  g1045
  (
    n992,
    n680
  );


  not
  g1046
  (
    n1033,
    n743
  );


  not
  g1047
  (
    n928,
    n692
  );


  buf
  g1048
  (
    n920,
    n643
  );


  not
  g1049
  (
    n862,
    n718
  );


  not
  g1050
  (
    n919,
    n670
  );


  buf
  g1051
  (
    n1070,
    n773
  );


  buf
  g1052
  (
    n970,
    n778
  );


  buf
  g1053
  (
    n1141,
    n882
  );


  not
  g1054
  (
    n1126,
    n863
  );


  not
  g1055
  (
    n1114,
    n884
  );


  not
  g1056
  (
    n1089,
    n865
  );


  not
  g1057
  (
    n1123,
    n890
  );


  buf
  g1058
  (
    n1121,
    n889
  );


  buf
  g1059
  (
    n1138,
    n910
  );


  buf
  g1060
  (
    n1115,
    n899
  );


  buf
  g1061
  (
    n1112,
    n886
  );


  not
  g1062
  (
    n1085,
    n866
  );


  buf
  g1063
  (
    n1087,
    n881
  );


  buf
  g1064
  (
    n1100,
    n862
  );


  buf
  g1065
  (
    n1097,
    n867
  );


  buf
  g1066
  (
    n1088,
    n902
  );


  not
  g1067
  (
    n1107,
    n893
  );


  not
  g1068
  (
    n1084,
    n909
  );


  buf
  g1069
  (
    n1124,
    n905
  );


  buf
  g1070
  (
    n1120,
    n912
  );


  buf
  g1071
  (
    n1113,
    n872
  );


  not
  g1072
  (
    n1118,
    n906
  );


  buf
  g1073
  (
    n1137,
    n868
  );


  buf
  g1074
  (
    n1117,
    n874
  );


  not
  g1075
  (
    n1140,
    n907
  );


  not
  g1076
  (
    n1106,
    n883
  );


  not
  g1077
  (
    n1131,
    n878
  );


  buf
  g1078
  (
    n1104,
    n880
  );


  buf
  g1079
  (
    n1092,
    n871
  );


  not
  g1080
  (
    n1091,
    n908
  );


  buf
  g1081
  (
    n1134,
    n876
  );


  not
  g1082
  (
    n1129,
    n903
  );


  buf
  g1083
  (
    n1127,
    n915
  );


  buf
  g1084
  (
    n1122,
    n894
  );


  not
  g1085
  (
    n1105,
    n873
  );


  not
  g1086
  (
    n1125,
    n896
  );


  not
  g1087
  (
    n1128,
    n877
  );


  not
  g1088
  (
    n1086,
    n891
  );


  buf
  g1089
  (
    n1103,
    n888
  );


  not
  g1090
  (
    n1108,
    n914
  );


  not
  g1091
  (
    n1109,
    n892
  );


  not
  g1092
  (
    n1102,
    n870
  );


  buf
  g1093
  (
    n1096,
    n911
  );


  not
  g1094
  (
    n1119,
    n879
  );


  buf
  g1095
  (
    n1132,
    n864
  );


  not
  g1096
  (
    n1099,
    n901
  );


  buf
  g1097
  (
    n1116,
    n860
  );


  buf
  g1098
  (
    n1135,
    n887
  );


  buf
  g1099
  (
    n1139,
    n869
  );


  buf
  g1100
  (
    n1095,
    n895
  );


  buf
  g1101
  (
    n1098,
    n898
  );


  buf
  g1102
  (
    n1090,
    n875
  );


  buf
  g1103
  (
    n1110,
    n861
  );


  buf
  g1104
  (
    n1094,
    n900
  );


  buf
  g1105
  (
    n1093,
    n897
  );


  not
  g1106
  (
    n1130,
    n904
  );


  buf
  g1107
  (
    n1136,
    n913
  );


  not
  g1108
  (
    n1101,
    n858
  );


  buf
  g1109
  (
    n1111,
    n859
  );


  buf
  g1110
  (
    n1133,
    n885
  );


  or
  g1111
  (
    n1164,
    n622,
    n620,
    n1105,
    n1098
  );


  nor
  g1112
  (
    n1147,
    n623,
    n625,
    n622,
    n929
  );


  nand
  g1113
  (
    n1149,
    n624,
    n918,
    n1093,
    n620
  );


  and
  g1114
  (
    n1148,
    n623,
    n622,
    n621
  );


  nand
  g1115
  (
    n1163,
    n1090,
    n1084,
    n627,
    n921
  );


  xnor
  g1116
  (
    n1144,
    n1094,
    n930,
    n1111,
    n1097
  );


  xor
  g1117
  (
    n1150,
    n925,
    n627,
    n618,
    n1091
  );


  and
  g1118
  (
    AntiSAT_key_wire,
    n623,
    n628,
    n927,
    n618
  );


  nor
  g1119
  (
    n1142,
    n934,
    n617,
    n1088,
    n931
  );


  nor
  g1120
  (
    n1151,
    n619,
    n621,
    n620,
    n624
  );


  or
  g1121
  (
    n1158,
    n624,
    n1100,
    n619,
    n1107
  );


  and
  g1122
  (
    n1161,
    n622,
    n1104,
    n1101,
    n939
  );


  nor
  g1123
  (
    n1153,
    n1103,
    n1109,
    n626,
    n1102
  );


  or
  g1124
  (
    n1159,
    n1092,
    n924,
    n937,
    n626
  );


  nand
  g1125
  (
    n1154,
    n627,
    n620,
    n617,
    n936
  );


  nor
  g1126
  (
    n1143,
    n1106,
    n916,
    n624,
    n1089
  );


  xnor
  g1127
  (
    n1165,
    n1086,
    n940,
    n621,
    n935
  );


  nor
  g1128
  (
    n1157,
    n628,
    n619,
    n618,
    n1110
  );


  xor
  g1129
  (
    n1160,
    n919,
    n628,
    n629,
    n920
  );


  xor
  g1130
  (
    n1166,
    n1085,
    n617,
    n933,
    n626
  );


  xor
  g1131
  (
    n1156,
    n629,
    n938,
    n917,
    n1096
  );


  xor
  g1132
  (
    n1146,
    n627,
    n626,
    n617,
    n1099
  );


  and
  g1133
  (
    n1162,
    n1095,
    n926,
    n1108,
    n928
  );


  nand
  g1134
  (
    n1145,
    n623,
    n923,
    n941,
    n625
  );


  and
  g1135
  (
    n1167,
    n625,
    n625,
    n618,
    n922
  );


  or
  g1136
  (
    n1155,
    n619,
    n932,
    n628,
    n1087
  );


  buf
  g1137
  (
    n1175,
    n1159
  );


  not
  g1138
  (
    n1173,
    n950
  );


  not
  g1139
  (
    n1168,
    n944
  );


  not
  g1140
  (
    n1170,
    n945
  );


  buf
  g1141
  (
    n1172,
    n1165
  );


  buf
  g1142
  (
    n1174,
    n948
  );


  not
  g1143
  (
    n1176,
    n1161
  );


  xor
  g1144
  (
    n1177,
    n1167,
    n1158,
    n947,
    n949
  );


  xnor
  g1145
  (
    n1169,
    n1164,
    n1163,
    n943,
    n1162
  );


  or
  g1146
  (
    n1171,
    n1160,
    n1166,
    n942,
    n946
  );


  nor
  g1147
  (
    n1182,
    n998,
    n1175,
    n1174,
    n980
  );


  xor
  g1148
  (
    n1193,
    n954,
    n1004,
    n991,
    n1175
  );


  nand
  g1149
  (
    n1186,
    n1175,
    n972,
    n968,
    n1002
  );


  nor
  g1150
  (
    n1181,
    n999,
    n958,
    n990,
    n993
  );


  nand
  g1151
  (
    n1188,
    n962,
    n973,
    n960,
    n1176
  );


  xnor
  g1152
  (
    n1183,
    n966,
    n981,
    n986,
    n995
  );


  or
  g1153
  (
    n1180,
    n1007,
    n965,
    n982,
    n956
  );


  or
  g1154
  (
    n1196,
    n1170,
    n1172,
    n1008,
    n996
  );


  xor
  g1155
  (
    n1179,
    n1174,
    n1171,
    n961,
    n976
  );


  or
  g1156
  (
    n1184,
    n1172,
    n1009,
    n957,
    n963
  );


  xor
  g1157
  (
    n1185,
    n952,
    n983,
    n974,
    n987
  );


  xnor
  g1158
  (
    n1191,
    n997,
    n1172,
    n1174,
    n994
  );


  or
  g1159
  (
    n1192,
    n1175,
    n989,
    n959,
    n979
  );


  xnor
  g1160
  (
    n1190,
    n988,
    n1174,
    n1003,
    n955
  );


  nor
  g1161
  (
    n1178,
    n978,
    n1173,
    n1176,
    n1000
  );


  and
  g1162
  (
    n1194,
    n1005,
    n1169,
    n1173,
    n1001
  );


  nor
  g1163
  (
    n1197,
    n984,
    n992,
    n969,
    n1010
  );


  xor
  g1164
  (
    n1195,
    n967,
    n970,
    n953,
    n971
  );


  xnor
  g1165
  (
    n1187,
    n985,
    n964,
    n951,
    n1006
  );


  xnor
  g1166
  (
    n1189,
    n975,
    n1168,
    n977,
    n1173
  );


  or
  g1167
  (
    n1202,
    n1021,
    n1023,
    n1113,
    n1122
  );


  xor
  g1168
  (
    n1208,
    n1184,
    n1115,
    n1116,
    n1122
  );


  xor
  g1169
  (
    n1199,
    n1022,
    n1187,
    n1115,
    n1116
  );


  xor
  g1170
  (
    n1209,
    n1195,
    n1189,
    n1118,
    n1122
  );


  nor
  g1171
  (
    n1201,
    n1118,
    n1124,
    n1114,
    n1119
  );


  nand
  g1172
  (
    n1198,
    n1019,
    n1119,
    n1013,
    n1121
  );


  nand
  g1173
  (
    n1200,
    n1117,
    n1119,
    n1118,
    n1121
  );


  xor
  g1174
  (
    n1207,
    n1114,
    n1120,
    n1012,
    n1191
  );


  or
  g1175
  (
    n1210,
    n1185,
    n1020,
    n1193,
    n1182
  );


  or
  g1176
  (
    n1213,
    n1117,
    n1015,
    n1186,
    n1120
  );


  nand
  g1177
  (
    n1206,
    n1011,
    n1197,
    n1014,
    n1114
  );


  nor
  g1178
  (
    n1205,
    n1024,
    n1194,
    n1120,
    n1018
  );


  xnor
  g1179
  (
    n1203,
    n1190,
    n1115,
    n1121,
    n1123
  );


  nand
  g1180
  (
    n1204,
    n1017,
    n1112,
    n1183,
    n1123
  );


  nand
  g1181
  (
    n1211,
    n1117,
    n1016,
    n1124,
    n1196
  );


  and
  g1182
  (
    n1212,
    n1123,
    n1116,
    n1188,
    n1192
  );


  not
  g1183
  (
    n1219,
    n1129
  );


  not
  g1184
  (
    n1224,
    n1133
  );


  not
  g1185
  (
    n1228,
    n1208
  );


  not
  g1186
  (
    n1222,
    n1199
  );


  or
  g1187
  (
    n1215,
    n1127,
    n1028,
    n1133
  );


  or
  g1188
  (
    n1225,
    n1128,
    n1129,
    n1126,
    n1201
  );


  xnor
  g1189
  (
    n1218,
    n1125,
    n1131,
    n1025,
    n1130
  );


  or
  g1190
  (
    n1214,
    n1132,
    n1128,
    n1205,
    n1207
  );


  xnor
  g1191
  (
    n1220,
    n1210,
    n1026,
    n1027,
    n1200
  );


  and
  g1192
  (
    n1226,
    n1204,
    n1212,
    n1198,
    n1130
  );


  xor
  g1193
  (
    n1227,
    n1202,
    n1127,
    n1206,
    n1125
  );


  nand
  g1194
  (
    n1221,
    n1130,
    n1132,
    n1209,
    n1127
  );


  and
  g1195
  (
    n1223,
    n1133,
    n1131,
    n1203,
    n1129
  );


  and
  g1196
  (
    n1216,
    n1124,
    n1126,
    n1125
  );


  or
  g1197
  (
    n1217,
    n1132,
    n1128,
    n1131,
    n1211
  );


  buf
  g1198
  (
    n1237,
    n1215
  );


  not
  g1199
  (
    n1243,
    n629
  );


  not
  g1200
  (
    n1240,
    n1228
  );


  not
  g1201
  (
    n1241,
    n1227
  );


  not
  g1202
  (
    n1235,
    n1214
  );


  not
  g1203
  (
    n1230,
    n630
  );


  not
  g1204
  (
    n1229,
    n1222
  );


  not
  g1205
  (
    n1233,
    n1217
  );


  not
  g1206
  (
    n1234,
    n630
  );


  not
  g1207
  (
    n1232,
    n629
  );


  not
  g1208
  (
    n1239,
    n1226
  );


  buf
  g1209
  (
    n1244,
    n1221
  );


  buf
  g1210
  (
    n1231,
    n1225
  );


  buf
  g1211
  (
    n1245,
    n1228
  );


  xnor
  g1212
  (
    n1238,
    n630,
    n1216
  );


  xor
  g1213
  (
    n1236,
    n1219,
    n1220,
    n1224
  );


  nand
  g1214
  (
    n1242,
    n1223,
    n1228,
    n1218
  );


  nor
  g1215
  (
    n1252,
    n1058,
    n1235
  );


  or
  g1216
  (
    n1247,
    n1030,
    n1245
  );


  xor
  g1217
  (
    n1272,
    n1042,
    n1240
  );


  and
  g1218
  (
    n1275,
    n1063,
    n1041
  );


  xor
  g1219
  (
    n1251,
    n1239,
    n1244
  );


  and
  g1220
  (
    n1274,
    n1239,
    n1232
  );


  nand
  g1221
  (
    n1258,
    n1241,
    n1230
  );


  and
  g1222
  (
    n1277,
    n1051,
    n1242
  );


  or
  g1223
  (
    n1280,
    n1055,
    n1245
  );


  xnor
  g1224
  (
    n1250,
    n1242,
    n1237
  );


  or
  g1225
  (
    n1278,
    n1031,
    n1243
  );


  nand
  g1226
  (
    n1249,
    n1243,
    n1035
  );


  or
  g1227
  (
    n1261,
    n1236,
    n1241
  );


  nor
  g1228
  (
    n1259,
    n1046,
    n1062
  );


  xnor
  g1229
  (
    n1246,
    n1029,
    n1245
  );


  nand
  g1230
  (
    n1267,
    n1060,
    n1240
  );


  and
  g1231
  (
    n1269,
    n1050,
    n857
  );


  and
  g1232
  (
    n1257,
    n1040,
    n1052
  );


  or
  g1233
  (
    n1279,
    n1243,
    n1241
  );


  or
  g1234
  (
    n1276,
    n1048,
    n1229
  );


  xor
  g1235
  (
    n1262,
    n1059,
    n1043
  );


  xnor
  g1236
  (
    n1270,
    n1233,
    n1241
  );


  and
  g1237
  (
    n1266,
    n1244,
    n1045
  );


  nor
  g1238
  (
    n1254,
    n1044,
    n1036
  );


  xnor
  g1239
  (
    n1260,
    n1034,
    n1054
  );


  nor
  g1240
  (
    n1255,
    n1244,
    n1056
  );


  nor
  g1241
  (
    n1268,
    n1049,
    n1239
  );


  or
  g1242
  (
    n1265,
    n1047,
    n1243
  );


  nor
  g1243
  (
    n1248,
    n1037,
    n1234
  );


  buf
  g1244
  (
    n1263,
    n1242
  );


  xor
  g1245
  (
    n1264,
    n1244,
    n1033
  );


  xor
  g1246
  (
    n1253,
    n1057,
    n1053
  );


  nand
  g1247
  (
    n1256,
    n1038,
    n1245
  );


  nand
  g1248
  (
    n1271,
    n1032,
    n1231
  );


  xnor
  g1249
  (
    n1281,
    n1039,
    n1240
  );


  or
  g1250
  (
    n1273,
    n1061,
    n1238
  );


  not
  g1251
  (
    n1283,
    n1261
  );


  not
  g1252
  (
    n1296,
    n1258
  );


  buf
  g1253
  (
    n1294,
    n1253
  );


  not
  g1254
  (
    n1290,
    n1252
  );


  buf
  g1255
  (
    n1297,
    n1249
  );


  buf
  g1256
  (
    n1291,
    n1250
  );


  not
  g1257
  (
    n1282,
    n1248
  );


  buf
  g1258
  (
    n1284,
    n1255
  );


  not
  g1259
  (
    n1295,
    n1257
  );


  buf
  g1260
  (
    n1286,
    n1247
  );


  not
  g1261
  (
    n1288,
    n1256
  );


  not
  g1262
  (
    n1287,
    n1254
  );


  buf
  g1263
  (
    n1289,
    n1251
  );


  buf
  g1264
  (
    n1293,
    n1260
  );


  not
  g1265
  (
    n1292,
    n1259
  );


  not
  g1266
  (
    n1285,
    n1246
  );


  not
  g1267
  (
    n1302,
    n1282
  );


  not
  g1268
  (
    n1298,
    n1133
  );


  nor
  g1269
  (
    n1300,
    n1282,
    n1065
  );


  nand
  g1270
  (
    n1303,
    n1283,
    n1066
  );


  nor
  g1271
  (
    n1301,
    n1064,
    n1282
  );


  xor
  g1272
  (
    n1299,
    n1283,
    n1282
  );


  xor
  g1273
  (
    n1305,
    n1299,
    n1072,
    n1074,
    n1298
  );


  nor
  g1274
  (
    n1304,
    n1134,
    n1301,
    n1070,
    n1068
  );


  nand
  g1275
  (
    n1307,
    n1300,
    n1073,
    n1067,
    n1071
  );


  nand
  g1276
  (
    n1306,
    n1069,
    n1134
  );


  xnor
  g1277
  (
    n1309,
    n1177,
    n1176,
    n1136
  );


  xor
  g1278
  (
    n1311,
    n1136,
    n1304,
    n1305
  );


  xnor
  g1279
  (
    n1310,
    n1137,
    n1076,
    n1177,
    n1136
  );


  xor
  g1280
  (
    n1308,
    n1305,
    n1304,
    n1135
  );


  xnor
  g1281
  (
    n1312,
    n1177,
    n1138,
    n1137,
    n1075
  );


  xor
  g1282
  (
    n1313,
    n1135,
    n1304,
    n1137
  );


  and
  g1283
  (
    n1314,
    n1177,
    n1136,
    n1305,
    n1135
  );


  and
  g1284
  (
    n1323,
    n1288,
    n1309
  );


  xnor
  g1285
  (
    n1328,
    n1289,
    n1286,
    n1312
  );


  and
  g1286
  (
    n1327,
    n1285,
    n1283,
    n1313
  );


  nor
  g1287
  (
    n1329,
    n1286,
    n1290,
    n1284
  );


  nand
  g1288
  (
    n1325,
    n1284,
    n1308,
    n1286
  );


  or
  g1289
  (
    n1316,
    n1314,
    n1288,
    n1289
  );


  nand
  g1290
  (
    n1319,
    n1310,
    n1314,
    n1285
  );


  and
  g1291
  (
    n1326,
    n1286,
    n1311,
    n1289
  );


  nand
  g1292
  (
    n1322,
    n1288,
    n1312,
    n1290
  );


  nand
  g1293
  (
    n1317,
    n1289,
    n1290,
    n1283
  );


  xnor
  g1294
  (
    n1320,
    n1313,
    n1287
  );


  and
  g1295
  (
    n1315,
    n1287,
    n1313
  );


  xor
  g1296
  (
    n1324,
    n1284,
    n1287,
    n1285
  );


  or
  g1297
  (
    n1318,
    n1312,
    n1288,
    n1284
  );


  nand
  g1298
  (
    n1321,
    n1285,
    n1314
  );


  xor
  g1299
  (
    n1344,
    n1324,
    n1141
  );


  xnor
  g1300
  (
    n1335,
    n1317,
    n1139
  );


  or
  g1301
  (
    n1342,
    n1321,
    n1329
  );


  xnor
  g1302
  (
    n1333,
    n1140,
    n1315,
    n1081
  );


  or
  g1303
  (
    n1338,
    n1290,
    n1323,
    n1329
  );


  or
  g1304
  (
    n1340,
    n1325,
    n1292,
    n1078
  );


  xor
  g1305
  (
    n1332,
    n1139,
    n1141,
    n1140
  );


  and
  g1306
  (
    n1339,
    n1291,
    n1322,
    n1079
  );


  nand
  g1307
  (
    n1334,
    n1327,
    n1291,
    n1328
  );


  nor
  g1308
  (
    n1337,
    n1082,
    n1139,
    n1316
  );


  nand
  g1309
  (
    n1331,
    n1292,
    n1303,
    n1139
  );


  xnor
  g1310
  (
    n1336,
    n1138,
    n1302,
    n1319
  );


  nor
  g1311
  (
    n1346,
    n1080,
    n1140,
    n1329
  );


  xor
  g1312
  (
    n1341,
    n1138,
    n1141
  );


  nand
  g1313
  (
    n1330,
    n1291,
    n1138,
    n1140
  );


  and
  g1314
  (
    n1345,
    n1292,
    n1320,
    n1077
  );


  nor
  g1315
  (
    n1343,
    n1291,
    n1318,
    n1326
  );


  buf
  g1316
  (
    n1357,
    n1273
  );


  not
  g1317
  (
    n1362,
    n1296
  );


  not
  g1318
  (
    n1360,
    n1265
  );


  buf
  g1319
  (
    n1351,
    n1295
  );


  xor
  g1320
  (
    n1359,
    n1296,
    n1333,
    n1271,
    n1346
  );


  xnor
  g1321
  (
    n1365,
    n1294,
    n1336,
    n1344,
    n1083
  );


  or
  g1322
  (
    n1364,
    n1339,
    n1266,
    n1269,
    n1296
  );


  or
  g1323
  (
    n1352,
    n1306,
    n1307,
    n1345
  );


  or
  g1324
  (
    n1355,
    n1306,
    n630,
    n1334,
    n1297
  );


  xnor
  g1325
  (
    n1349,
    n1294,
    n1264,
    n1346,
    n1341
  );


  xnor
  g1326
  (
    n1348,
    n1295,
    n1293,
    n1346,
    n1332
  );


  or
  g1327
  (
    n1350,
    n1268,
    n1337,
    n1306,
    n1213
  );


  or
  g1328
  (
    n1354,
    n1342,
    n1294,
    n1330,
    n1295
  );


  xnor
  g1329
  (
    n1358,
    n1297,
    n1338,
    n1263,
    n1292
  );


  or
  g1330
  (
    n1356,
    n1272,
    n1307,
    n1294,
    n1297
  );


  xor
  g1331
  (
    n1363,
    n1340,
    n1293,
    n1267
  );


  xor
  g1332
  (
    n1361,
    n1293,
    n1331,
    n1295,
    n1297
  );


  xor
  g1333
  (
    n1347,
    n1306,
    n1270,
    n1343,
    n1296
  );


  nor
  g1334
  (
    n1353,
    n1307,
    n1305,
    n1335,
    n1262
  );


  not
  g1335
  (
    n1383,
    n1356
  );


  buf
  g1336
  (
    n1439,
    n1364
  );


  not
  g1337
  (
    n1438,
    n1349
  );


  not
  g1338
  (
    n1401,
    n1352
  );


  buf
  g1339
  (
    n1375,
    n1353
  );


  buf
  g1340
  (
    n1433,
    n1364
  );


  buf
  g1341
  (
    n1404,
    n1349
  );


  not
  g1342
  (
    n1395,
    n1365
  );


  not
  g1343
  (
    n1379,
    n1351
  );


  not
  g1344
  (
    n1434,
    n1360
  );


  buf
  g1345
  (
    n1377,
    n1349
  );


  not
  g1346
  (
    n1373,
    n1360
  );


  not
  g1347
  (
    n1426,
    n1350
  );


  not
  g1348
  (
    n1407,
    n1363
  );


  not
  g1349
  (
    n1409,
    n1364
  );


  not
  g1350
  (
    n1431,
    n1359
  );


  not
  g1351
  (
    n1386,
    n1361
  );


  buf
  g1352
  (
    n1382,
    n1348
  );


  not
  g1353
  (
    n1435,
    n1358
  );


  buf
  g1354
  (
    n1425,
    n1356
  );


  buf
  g1355
  (
    n1372,
    n1355
  );


  buf
  g1356
  (
    n1392,
    n1360
  );


  buf
  g1357
  (
    n1393,
    n1352
  );


  buf
  g1358
  (
    n1400,
    n1351
  );


  not
  g1359
  (
    n1410,
    n1354
  );


  buf
  g1360
  (
    n1405,
    n1351
  );


  buf
  g1361
  (
    n1391,
    n1354
  );


  not
  g1362
  (
    n1368,
    n1358
  );


  buf
  g1363
  (
    n1378,
    n1352
  );


  not
  g1364
  (
    n1419,
    n1362
  );


  not
  g1365
  (
    n1441,
    n1365
  );


  not
  g1366
  (
    n1389,
    n1361
  );


  buf
  g1367
  (
    n1396,
    n1347
  );


  not
  g1368
  (
    n1436,
    n1353
  );


  not
  g1369
  (
    n1398,
    n1362
  );


  buf
  g1370
  (
    n1369,
    n1347
  );


  not
  g1371
  (
    n1406,
    n1360
  );


  not
  g1372
  (
    n1370,
    n1354
  );


  not
  g1373
  (
    n1390,
    n1358
  );


  buf
  g1374
  (
    n1416,
    n1357
  );


  buf
  g1375
  (
    n1424,
    n1347
  );


  buf
  g1376
  (
    n1380,
    n1359
  );


  not
  g1377
  (
    n1376,
    n1357
  );


  buf
  g1378
  (
    n1414,
    n1355
  );


  buf
  g1379
  (
    n1428,
    n1350
  );


  not
  g1380
  (
    n1374,
    n1355
  );


  not
  g1381
  (
    n1387,
    n1365
  );


  buf
  g1382
  (
    n1412,
    n1350
  );


  buf
  g1383
  (
    n1394,
    n1359
  );


  buf
  g1384
  (
    n1440,
    n1363
  );


  buf
  g1385
  (
    n1437,
    n1348
  );


  buf
  g1386
  (
    n1367,
    n1363
  );


  not
  g1387
  (
    n1421,
    n1364
  );


  buf
  g1388
  (
    n1427,
    n1362
  );


  not
  g1389
  (
    n1418,
    n1357
  );


  buf
  g1390
  (
    n1411,
    n1359
  );


  buf
  g1391
  (
    n1429,
    n1352
  );


  buf
  g1392
  (
    n1422,
    n1348
  );


  not
  g1393
  (
    n1408,
    n1356
  );


  buf
  g1394
  (
    n1385,
    n1356
  );


  not
  g1395
  (
    n1397,
    n1355
  );


  not
  g1396
  (
    n1420,
    n1361
  );


  not
  g1397
  (
    n1403,
    n1353
  );


  buf
  g1398
  (
    n1402,
    n1357
  );


  not
  g1399
  (
    n1388,
    n1361
  );


  not
  g1400
  (
    n1366,
    n1353
  );


  not
  g1401
  (
    n1417,
    n1347
  );


  not
  g1402
  (
    n1415,
    n1358
  );


  not
  g1403
  (
    n1413,
    n1351
  );


  buf
  g1404
  (
    n1384,
    n1365
  );


  buf
  g1405
  (
    n1423,
    n1363
  );


  not
  g1406
  (
    n1430,
    n1354
  );


  not
  g1407
  (
    n1432,
    n1362
  );


  not
  g1408
  (
    n1371,
    n1350
  );


  not
  g1409
  (
    n1381,
    n1349
  );


  not
  g1410
  (
    n1399,
    n1348
  );


  and
  g1411
  (
    n1455,
    n1439,
    n1368,
    n1437,
    n1279
  );


  nor
  g1412
  (
    n1449,
    n1407,
    n1420,
    n1279
  );


  or
  g1413
  (
    n1462,
    n1369,
    n1437,
    n1439,
    n1395
  );


  or
  g1414
  (
    n1444,
    n1434,
    n1427,
    n1417,
    n1422
  );


  or
  g1415
  (
    n1446,
    n1401,
    n1387,
    n1439,
    n1419
  );


  and
  g1416
  (
    n1453,
    n1280,
    n1423,
    n1406,
    n1432
  );


  nor
  g1417
  (
    n1469,
    n1438,
    n1441,
    n1373,
    n1430
  );


  xnor
  g1418
  (
    n1442,
    n1386,
    n1425,
    n1410,
    n1428
  );


  or
  g1419
  (
    n1465,
    n1391,
    n1438,
    n1366,
    n1378
  );


  xnor
  g1420
  (
    n1473,
    n1276,
    n1398,
    n1388,
    n1433
  );


  nor
  g1421
  (
    n1468,
    n1416,
    n1278,
    n1432,
    n1400
  );


  nand
  g1422
  (
    n1452,
    n1429,
    n1276,
    n1379,
    n1435
  );


  and
  g1423
  (
    n1451,
    n1415,
    n1372,
    n1433,
    n1426
  );


  and
  g1424
  (
    n1459,
    n1377,
    n1280,
    n1279,
    n1434
  );


  xor
  g1425
  (
    n1475,
    n1422,
    n1428,
    n1367,
    n1421
  );


  and
  g1426
  (
    n1467,
    n1374,
    n1426,
    n1425,
    n1275
  );


  and
  g1427
  (
    n1461,
    n1279,
    n1402,
    n1435,
    n1441
  );


  and
  g1428
  (
    n1471,
    n1423,
    n1434,
    n1431,
    n1381
  );


  nor
  g1429
  (
    n1448,
    n1413,
    n1418,
    n1276,
    n1280
  );


  or
  g1430
  (
    n1443,
    n1277,
    n1370,
    n1394,
    n1436
  );


  or
  g1431
  (
    n1450,
    n1382,
    n1281,
    n1431,
    n1420
  );


  nor
  g1432
  (
    n1470,
    n1384,
    n1405,
    n1277,
    n1414
  );


  or
  g1433
  (
    n1456,
    n1436,
    n1433,
    n1380,
    n1424
  );


  nor
  g1434
  (
    n1476,
    n1278,
    n1440,
    n1383,
    n1376
  );


  xor
  g1435
  (
    n1463,
    n1427,
    n1430,
    n1392,
    n1425
  );


  or
  g1436
  (
    n1454,
    n1385,
    n1397,
    n1277,
    n1440
  );


  xnor
  g1437
  (
    n1447,
    n1399,
    n1390,
    n1409,
    n1278
  );


  xor
  g1438
  (
    n1460,
    n1436,
    n1396,
    n1435,
    n1423
  );


  xnor
  g1439
  (
    n1477,
    n1426,
    n1403,
    n1411,
    n1281
  );


  and
  g1440
  (
    n1474,
    n1432,
    n1389,
    n1404,
    n1281
  );


  xor
  g1441
  (
    n1472,
    n1393,
    n1431,
    n1429,
    n1281
  );


  nor
  g1442
  (
    n1445,
    n1375,
    n1437,
    n1421,
    n1424
  );


  xor
  g1443
  (
    n1464,
    n1441,
    n1371,
    n1427,
    n1438
  );


  or
  g1444
  (
    n1457,
    n1280,
    n1430,
    n1274,
    n1424
  );


  xnor
  g1445
  (
    n1466,
    n1440,
    n1429,
    n1422,
    n1428
  );


  and
  g1446
  (
    n1458,
    n1408,
    n1421,
    n1278,
    n1412
  );


  nand
  g1447
  (
    n1481,
    n1443,
    n1471,
    n1477,
    n1470
  );


  xnor
  g1448
  (
    n1486,
    n1465,
    n1472,
    n1457,
    n1448
  );


  nor
  g1449
  (
    n1484,
    n1461,
    n1467,
    n1466,
    n1452
  );


  nand
  g1450
  (
    n1480,
    n1463,
    n1456,
    n1451,
    n1455
  );


  xnor
  g1451
  (
    n1485,
    n1446,
    n1473,
    n1458,
    n1449
  );


  xnor
  g1452
  (
    n1479,
    n1447,
    n1442,
    n1469,
    n1474
  );


  or
  g1453
  (
    n1483,
    n1475,
    n1453,
    n1445,
    n1460
  );


  xnor
  g1454
  (
    n1478,
    n1454,
    n1450,
    n1444,
    n1468
  );


  xnor
  g1455
  (
    n1482,
    n1464,
    n1476,
    n1462,
    n1459
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_30
  (
    gbar_input_0_0,
    keyIn_0_30,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_1,
    keyIn_0_31,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_2,
    keyIn_0_32,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_3,
    keyIn_0_33,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_4,
    keyIn_0_34,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_5,
    keyIn_0_35,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_6,
    keyIn_0_36,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_7,
    keyIn_0_37,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_8,
    keyIn_0_38,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_9,
    keyIn_0_39,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_10,
    keyIn_0_40,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_11,
    keyIn_0_41,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_12,
    keyIn_0_42,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_13,
    keyIn_0_43,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_14,
    keyIn_0_44,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_15,
    keyIn_0_45,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_16,
    keyIn_0_46,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_17,
    keyIn_0_47,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_18,
    keyIn_0_48,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_19,
    keyIn_0_49,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_20,
    keyIn_0_50,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_21,
    keyIn_0_51,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_22,
    keyIn_0_52,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_23,
    keyIn_0_53,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_24,
    keyIn_0_54,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_25,
    keyIn_0_55,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_26,
    keyIn_0_56,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_27,
    keyIn_0_57,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_28,
    keyIn_0_58,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_29,
    keyIn_0_59,
    n30
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n1152,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

