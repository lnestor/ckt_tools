// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_58 written by SynthGen on 2021/04/05 11:22:31
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_58 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n112, n108, n113, n110, n105, n128, n129, n131,
 n107, n122, n118, n115, n127, n130, n121, n102,
 n103, n106, n132, n124, n104, n125, n119, n123,
 n116, n117, n120, n109, n126, n101, n114, n111);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n112, n108, n113, n110, n105, n128, n129, n131,
 n107, n122, n118, n115, n127, n130, n121, n102,
 n103, n106, n132, n124, n104, n125, n119, n123,
 n116, n117, n120, n109, n126, n101, n114, n111;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100;

buf  g0 (n63, n17);
not  g1 (n53, n16);
buf  g2 (n70, n13);
not  g3 (n45, n13);
buf  g4 (n66, n10);
not  g5 (n49, n12);
not  g6 (n67, n16);
buf  g7 (n58, n9);
not  g8 (n46, n15);
buf  g9 (n42, n17);
buf  g10 (n61, n14);
buf  g11 (n50, n18);
buf  g12 (n71, n1);
not  g13 (n40, n14);
buf  g14 (n72, n18);
not  g15 (n43, n5);
buf  g16 (n55, n19);
not  g17 (n48, n17);
not  g18 (n52, n11);
not  g19 (n65, n16);
buf  g20 (n47, n9);
not  g21 (n62, n11);
not  g22 (n41, n8);
not  g23 (n56, n11);
buf  g24 (n39, n4);
buf  g25 (n35, n12);
not  g26 (n38, n3);
not  g27 (n36, n12);
buf  g28 (n34, n19);
buf  g29 (n57, n6);
buf  g30 (n68, n9);
not  g31 (n37, n13);
buf  g32 (n69, n18);
buf  g33 (n44, n2);
buf  g34 (n33, n7);
not  g35 (n64, n15);
buf  g36 (n59, n15);
not  g37 (n51, n10);
buf  g38 (n54, n14);
buf  g39 (n60, n10);
buf  g40 (n77, n37);
buf  g41 (n76, n40);
buf  g42 (n80, n38);
buf  g43 (n78, n34);
not  g44 (n75, n36);
buf  g45 (n74, n40);
not  g46 (n79, n35);
nor  g47 (n73, n33, n39, n40);
buf  g48 (n82, n73);
not  g49 (n84, n75);
not  g50 (n83, n74);
not  g51 (n85, n77);
not  g52 (n81, n76);
nand g53 (n96, n22, n80, n81, n27);
and  g54 (n98, n32, n21, n84);
xnor g55 (n91, n24, n78, n27, n20);
xnor g56 (n99, n30, n85, n32);
nand g57 (n88, n19, n25, n84, n24);
nor  g58 (n97, n22, n84, n32, n21);
xnor g59 (n100, n85, n29, n23, n82);
xor  g60 (n93, n80, n83, n31, n81);
xor  g61 (n94, n82, n31, n27);
xor  g62 (n86, n22, n25, n83, n26);
nand g63 (n87, n30, n30, n25, n20);
and  g64 (n89, n23, n26, n83, n82);
and  g65 (n90, n20, n79, n28, n29);
nor  g66 (n95, n23, n26, n29, n24);
or   g67 (n92, n81, n28, n80);
nor  g68 (n121, n44, n65, n56, n63);
and  g69 (n108, n59, n52, n45, n72);
xor  g70 (n126, n67, n62, n86, n98);
and  g71 (n123, n49, n59, n65, n55);
or   g72 (n109, n93, n69, n96);
nand g73 (n132, n54, n70, n92, n58);
xor  g74 (n106, n69, n43, n94, n62);
and  g75 (n125, n95, n61, n93, n42);
xor  g76 (n129, n53, n59, n60, n54);
or   g77 (n130, n94, n51, n64, n66);
nand g78 (n124, n46, n57, n92, n47);
xnor g79 (n119, n93, n72, n98, n71);
or   g80 (n107, n56, n97, n50, n64);
nor  g81 (n122, n42, n55, n53, n63);
and  g82 (n116, n52, n100, n97, n91);
nor  g83 (n114, n99, n94, n100, n57);
nor  g84 (n110, n98, n45, n69, n61);
or   g85 (n102, n95, n70, n87, n68);
xor  g86 (n111, n50, n49, n43, n71);
and  g87 (n104, n48, n56, n67, n51);
or   g88 (n131, n61, n41, n90, n70);
xnor g89 (n118, n48, n62, n64, n57);
and  g90 (n113, n50, n51, n44, n41);
xor  g91 (n120, n45, n66, n49, n99);
nand g92 (n105, n60, n52, n42, n97);
nand g93 (n115, n96, n68, n65, n63);
and  g94 (n112, n71, n67, n89, n53);
nor  g95 (n128, n66, n72, n55, n100);
or   g96 (n117, n46, n68, n43, n47);
or   g97 (n101, n58, n41, n95, n54);
nand g98 (n127, n44, n88, n58, n60);
nor  g99 (n103, n48, n99, n47, n46);
endmodule
