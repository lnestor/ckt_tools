module MyNand(a, b, c);
input b, c;
output a;
Nand NAND2(a, b, c);
endmodule

module MyNand3(a, b, c, d);
input b, c, d;
output a;
Nand NAND3(a, b, c, d);
endmodule

module MyNand4(a, b, c, d, e);
input b, c, d, e;
output a;
Nand NAND4(a, b, c, d, e);
endmodule

module MyNand8(a, b, c, d, e, f, g, h, i);
input b, c, d, e, f, g, h, i;
output a;
Nand NAND8(a, b, c, d, e, f, g, h, i);
endmodule

module MyNand5(a, b, c, d, e, f);
input b, c, d, e, f;
output a;
Nand NAND5(a, b, c, d, e, f);
endmodule

module MyAnd(a, b, c);
input b, c;
output a;
And AND2(a, b, c);
endmodule

module MyAnd3(a, b, c, d);
input b, c, d;
output a;
And AND3(a, b, c, d);
endmodule

module MyAnd4(a, b, c, d, e);
input b, c, d, e;
output a;
And AND4(a, b, c, d, e);
endmodule

module MyAnd5(a, b, c, d, e, f);
input b, c, d, e, f;
output a;
And AND5(a, b, c, d, e, f);
endmodule

module MyAnd8(a, b, c, d, e, f, g, h, i);
input b, c, d, e, f, g, h, i;
output a;
And AND8(a, b, c, d, e, f, g, h, i);
endmodule

module MyNor(a, b, c);
input b, c;
output a;
Nor NOR1(a, b, c);
endmodule

module MyBuf(a, b);
input b;
output a;
Buf BUF1(a, b);
endmodule

module MyNot(a, b);
input b;
output a;
Not NOT1(a, b);
endmodule

module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;

output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898;

MyNot NOT1_1 (N190, N1);
MyNot NOT1_2 (N194, N4);
MyNot NOT1_3 (N197, N7);
MyNot NOT1_4 (N201, N10);
MyNot NOT1_5 (N206, N13);
MyNot NOT1_6 (N209, N16);
MyNot NOT1_7 (N212, N19);
MyNot NOT1_8 (N216, N22);
MyNot NOT1_9 (N220, N25);
MyNot NOT1_10 (N225, N28);
MyNot NOT1_11 (N229, N31);
MyNot NOT1_12 (N232, N34);
MyNot NOT1_13 (N235, N37);
MyNot NOT1_14 (N239, N40);
MyNot NOT1_15 (N243, N43);
MyNot NOT1_16 (N247, N46);
MyNand NAND2_17 (N251, N63, N88);
MyNand NAND2_18 (N252, N66, N91);
MyNot NOT1_19 (N253, N72);
MyNot NOT1_20 (N256, N72);
MyBuf BUFF1_21 (N257, N69);
MyBuf BUFF1_22 (N260, N69);
MyNot NOT1_23 (N263, N76);
MyNot NOT1_24 (N266, N79);
MyNot NOT1_25 (N269, N82);
MyNot NOT1_26 (N272, N85);
MyNot NOT1_27 (N275, N104);
MyNot NOT1_28 (N276, N104);
MyNot NOT1_29 (N277, N88);
MyNot NOT1_30 (N280, N91);
MyBuf BUFF1_31 (N283, N94);
MyNot NOT1_32 (N290, N94);
MyBuf BUFF1_33 (N297, N94);
MyNot NOT1_34 (N300, N94);
MyBuf BUFF1_35 (N303, N99);
MyNot NOT1_36 (N306, N99);
MyNot NOT1_37 (N313, N99);
MyBuf BUFF1_38 (N316, N104);
MyNot NOT1_39 (N319, N104);
MyBuf BUFF1_40 (N326, N104);
MyBuf BUFF1_41 (N331, N104);
MyNot NOT1_42 (N338, N104);
MyBuf BUFF1_43 (N343, N1);
MyBuf BUFF1_44 (N346, N4);
MyBuf BUFF1_45 (N349, N7);
MyBuf BUFF1_46 (N352, N10);
MyBuf BUFF1_47 (N355, N13);
MyBuf BUFF1_48 (N358, N16);
MyBuf BUFF1_49 (N361, N19);
MyBuf BUFF1_50 (N364, N22);
MyBuf BUFF1_51 (N367, N25);
MyBuf BUFF1_52 (N370, N28);
MyBuf BUFF1_53 (N373, N31);
MyBuf BUFF1_54 (N376, N34);
MyBuf BUFF1_55 (N379, N37);
MyBuf BUFF1_56 (N382, N40);
MyBuf BUFF1_57 (N385, N43);
MyBuf BUFF1_58 (N388, N46);
MyNot NOT1_59 (N534, N343);
MyNot NOT1_60 (N535, N346);
MyNot NOT1_61 (N536, N349);
MyNot NOT1_62 (N537, N352);
MyNot NOT1_63 (N538, N355);
MyNot NOT1_64 (N539, N358);
MyNot NOT1_65 (N540, N361);
MyNot NOT1_66 (N541, N364);
MyNot NOT1_67 (N542, N367);
MyNot NOT1_68 (N543, N370);
MyNot NOT1_69 (N544, N373);
MyNot NOT1_70 (N545, N376);
MyNot NOT1_71 (N546, N379);
MyNot NOT1_72 (N547, N382);
MyNot NOT1_73 (N548, N385);
MyNot NOT1_74 (N549, N388);
MyNand NAND2_75 (N550, N306, N331);
MyNand NAND2_76 (N551, N306, N331);
MyNand NAND2_77 (N552, N306, N331);
MyNand NAND2_78 (N553, N306, N331);
MyNand NAND2_79 (N554, N306, N331);
MyNand NAND2_80 (N555, N306, N331);
MyBuf BUFF1_81 (N556, N190);
MyBuf BUFF1_82 (N559, N194);
MyBuf BUFF1_83 (N562, N206);
MyBuf BUFF1_84 (N565, N209);
MyBuf BUFF1_85 (N568, N225);
MyBuf BUFF1_86 (N571, N243);
MyAnd AND2_87 (N574, N63, N319);
MyBuf BUFF1_88 (N577, N220);
MyBuf BUFF1_89 (N580, N229);
MyBuf BUFF1_90 (N583, N232);
MyAnd AND2_91 (N586, N66, N319);
MyBuf BUFF1_92 (N589, N239);
MyAnd3 AND3_93 (N592, N49, N253, N319);
MyBuf BUFF1_94 (N595, N247);
MyBuf BUFF1_95 (N598, N239);
MyNand NAND2_96 (N601, N326, N277);
MyNand NAND2_97 (N602, N326, N280);
MyNand NAND2_98 (N603, N260, N72);
MyNand NAND2_99 (N608, N260, N300);
MyNand NAND2_100 (N612, N256, N300);
MyBuf BUFF1_101 (N616, N201);
MyBuf BUFF1_102 (N619, N216);
MyBuf BUFF1_103 (N622, N220);
MyBuf BUFF1_104 (N625, N239);
MyBuf BUFF1_105 (N628, N190);
MyBuf BUFF1_106 (N631, N190);
MyBuf BUFF1_107 (N634, N194);
MyBuf BUFF1_108 (N637, N229);
MyBuf BUFF1_109 (N640, N197);
MyAnd3 AND3_110 (N643, N56, N257, N319);
MyBuf BUFF1_111 (N646, N232);
MyBuf BUFF1_112 (N649, N201);
MyBuf BUFF1_113 (N652, N235);
MyAnd3 AND3_114 (N655, N60, N257, N319);
MyBuf BUFF1_115 (N658, N263);
MyBuf BUFF1_116 (N661, N263);
MyBuf BUFF1_117 (N664, N266);
MyBuf BUFF1_118 (N667, N266);
MyBuf BUFF1_119 (N670, N269);
MyBuf BUFF1_120 (N673, N269);
MyBuf BUFF1_121 (N676, N272);
MyBuf BUFF1_122 (N679, N272);
MyAnd AND2_123 (N682, N251, N316);
MyAnd AND2_124 (N685, N252, N316);
MyBuf BUFF1_125 (N688, N197);
MyBuf BUFF1_126 (N691, N197);
MyBuf BUFF1_127 (N694, N212);
MyBuf BUFF1_128 (N697, N212);
MyBuf BUFF1_129 (N700, N247);
MyBuf BUFF1_130 (N703, N247);
MyBuf BUFF1_131 (N706, N235);
MyBuf BUFF1_132 (N709, N235);
MyBuf BUFF1_133 (N712, N201);
MyBuf BUFF1_134 (N715, N201);
MyBuf BUFF1_135 (N718, N206);
MyBuf BUFF1_136 (N721, N216);
MyAnd3 AND3_137 (N724, N53, N253, N319);
MyBuf BUFF1_138 (N727, N243);
MyBuf BUFF1_139 (N730, N220);
MyBuf BUFF1_140 (N733, N220);
MyBuf BUFF1_141 (N736, N209);
MyBuf BUFF1_142 (N739, N216);
MyBuf BUFF1_143 (N742, N225);
MyBuf BUFF1_144 (N745, N243);
MyBuf BUFF1_145 (N748, N212);
MyBuf BUFF1_146 (N751, N225);
MyNot NOT1_147 (N886, N682);
MyNot NOT1_148 (N887, N685);
MyNot NOT1_149 (N888, N616);
MyNot NOT1_150 (N889, N619);
MyNot NOT1_151 (N890, N622);
MyNot NOT1_152 (N891, N625);
MyNot NOT1_153 (N892, N631);
MyNot NOT1_154 (N893, N643);
MyNot NOT1_155 (N894, N649);
MyNot NOT1_156 (N895, N652);
MyNot NOT1_157 (N896, N655);
MyAnd AND2_158 (N897, N49, N612);
MyAnd AND2_159 (N898, N56, N608);
MyNand NAND2_160 (N899, N53, N612);
MyNand NAND2_161 (N903, N60, N608);
MyNand NAND2_162 (N907, N49, N612);
MyNand NAND2_163 (N910, N56, N608);
MyNot NOT1_164 (N913, N661);
MyNot NOT1_165 (N914, N658);
MyNot NOT1_166 (N915, N667);
MyNot NOT1_167 (N916, N664);
MyNot NOT1_168 (N917, N673);
MyNot NOT1_169 (N918, N670);
MyNot NOT1_170 (N919, N679);
MyNot NOT1_171 (N920, N676);
MyNand4 NAND4_172 (N921, N277, N297, N326, N603);
MyNand4 NAND4_173 (N922, N280, N297, N326, N603);
MyNand3 NAND3_174 (N923, N303, N338, N603);
MyAnd3 AND3_175 (N926, N303, N338, N603);
MyBuf BUFF1_176 (N935, N556);
MyNot NOT1_177 (N938, N688);
MyBuf BUFF1_178 (N939, N556);
MyNot NOT1_179 (N942, N691);
MyBuf BUFF1_180 (N943, N562);
MyNot NOT1_181 (N946, N694);
MyBuf BUFF1_182 (N947, N562);
MyNot NOT1_183 (N950, N697);
MyBuf BUFF1_184 (N951, N568);
MyNot NOT1_185 (N954, N700);
MyBuf BUFF1_186 (N955, N568);
MyNot NOT1_187 (N958, N703);
MyBuf BUFF1_188 (N959, N574);
MyBuf BUFF1_189 (N962, N574);
MyBuf BUFF1_190 (N965, N580);
MyNot NOT1_191 (N968, N706);
MyBuf BUFF1_192 (N969, N580);
MyNot NOT1_193 (N972, N709);
MyBuf BUFF1_194 (N973, N586);
MyNot NOT1_195 (N976, N712);
MyBuf BUFF1_196 (N977, N586);
MyNot NOT1_197 (N980, N715);
MyBuf BUFF1_198 (N981, N592);
MyNot NOT1_199 (N984, N628);
MyBuf BUFF1_200 (N985, N592);
MyNot NOT1_201 (N988, N718);
MyNot NOT1_202 (N989, N721);
MyNot NOT1_203 (N990, N634);
MyNot NOT1_204 (N991, N724);
MyNot NOT1_205 (N992, N727);
MyNot NOT1_206 (N993, N637);
MyBuf BUFF1_207 (N994, N595);
MyNot NOT1_208 (N997, N730);
MyBuf BUFF1_209 (N998, N595);
MyNot NOT1_210 (N1001, N733);
MyNot NOT1_211 (N1002, N736);
MyNot NOT1_212 (N1003, N739);
MyNot NOT1_213 (N1004, N640);
MyNot NOT1_214 (N1005, N742);
MyNot NOT1_215 (N1006, N745);
MyNot NOT1_216 (N1007, N646);
MyNot NOT1_217 (N1008, N748);
MyNot NOT1_218 (N1009, N751);
MyBuf BUFF1_219 (N1010, N559);
MyBuf BUFF1_220 (N1013, N559);
MyBuf BUFF1_221 (N1016, N565);
MyBuf BUFF1_222 (N1019, N565);
MyBuf BUFF1_223 (N1022, N571);
MyBuf BUFF1_224 (N1025, N571);
MyBuf BUFF1_225 (N1028, N577);
MyBuf BUFF1_226 (N1031, N577);
MyBuf BUFF1_227 (N1034, N583);
MyBuf BUFF1_228 (N1037, N583);
MyBuf BUFF1_229 (N1040, N589);
MyBuf BUFF1_230 (N1043, N589);
MyBuf BUFF1_231 (N1046, N598);
MyBuf BUFF1_232 (N1049, N598);
MyNand NAND2_233 (N1054, N619, N888);
MyNand NAND2_234 (N1055, N616, N889);
MyNand NAND2_235 (N1063, N625, N890);
MyNand NAND2_236 (N1064, N622, N891);
MyNand NAND2_237 (N1067, N655, N895);
MyNand NAND2_238 (N1068, N652, N896);
MyNand NAND2_239 (N1119, N721, N988);
MyNand NAND2_240 (N1120, N718, N989);
MyNand NAND2_241 (N1121, N727, N991);
MyNand NAND2_242 (N1122, N724, N992);
MyNand NAND2_243 (N1128, N739, N1002);
MyNand NAND2_244 (N1129, N736, N1003);
MyNand NAND2_245 (N1130, N745, N1005);
MyNand NAND2_246 (N1131, N742, N1006);
MyNand NAND2_247 (N1132, N751, N1008);
MyNand NAND2_248 (N1133, N748, N1009);
MyNot NOT1_249 (N1148, N939);
MyNot NOT1_250 (N1149, N935);
MyNand NAND2_251 (N1150, N1054, N1055);
MyNot NOT1_252 (N1151, N943);
MyNot NOT1_253 (N1152, N947);
MyNot NOT1_254 (N1153, N955);
MyNot NOT1_255 (N1154, N951);
MyNot NOT1_256 (N1155, N962);
MyNot NOT1_257 (N1156, N969);
MyNot NOT1_258 (N1157, N977);
MyNand NAND2_259 (N1158, N1063, N1064);
MyNot NOT1_260 (N1159, N985);
MyNand NAND2_261 (N1160, N985, N892);
MyNot NOT1_262 (N1161, N998);
MyNand NAND2_263 (N1162, N1067, N1068);
MyNot NOT1_264 (N1163, N899);
MyBuf BUFF1_265 (N1164, N899);
MyNot NOT1_266 (N1167, N903);
MyBuf BUFF1_267 (N1168, N903);
MyNand NAND2_268 (N1171, N921, N923);
MyNand NAND2_269 (N1188, N922, N923);
MyNot NOT1_270 (N1205, N1010);
MyNand NAND2_271 (N1206, N1010, N938);
MyNot NOT1_272 (N1207, N1013);
MyNand NAND2_273 (N1208, N1013, N942);
MyNot NOT1_274 (N1209, N1016);
MyNand NAND2_275 (N1210, N1016, N946);
MyNot NOT1_276 (N1211, N1019);
MyNand NAND2_277 (N1212, N1019, N950);
MyNot NOT1_278 (N1213, N1022);
MyNand NAND2_279 (N1214, N1022, N954);
MyNot NOT1_280 (N1215, N1025);
MyNand NAND2_281 (N1216, N1025, N958);
MyNot NOT1_282 (N1217, N1028);
MyNot NOT1_283 (N1218, N959);
MyNot NOT1_284 (N1219, N1031);
MyNot NOT1_285 (N1220, N1034);
MyNand NAND2_286 (N1221, N1034, N968);
MyNot NOT1_287 (N1222, N965);
MyNot NOT1_288 (N1223, N1037);
MyNand NAND2_289 (N1224, N1037, N972);
MyNot NOT1_290 (N1225, N1040);
MyNand NAND2_291 (N1226, N1040, N976);
MyNot NOT1_292 (N1227, N973);
MyNot NOT1_293 (N1228, N1043);
MyNand NAND2_294 (N1229, N1043, N980);
MyNot NOT1_295 (N1230, N981);
MyNand NAND2_296 (N1231, N981, N984);
MyNand NAND2_297 (N1232, N1119, N1120);
MyNand NAND2_298 (N1235, N1121, N1122);
MyNot NOT1_299 (N1238, N1046);
MyNand NAND2_300 (N1239, N1046, N997);
MyNot NOT1_301 (N1240, N994);
MyNot NOT1_302 (N1241, N1049);
MyNand NAND2_303 (N1242, N1049, N1001);
MyNand NAND2_304 (N1243, N1128, N1129);
MyNand NAND2_305 (N1246, N1130, N1131);
MyNand NAND2_306 (N1249, N1132, N1133);
MyBuf BUFF1_307 (N1252, N907);
MyBuf BUFF1_308 (N1255, N907);
MyBuf BUFF1_309 (N1258, N910);
MyBuf BUFF1_310 (N1261, N910);
MyNot NOT1_311 (N1264, N1150);
MyNand NAND2_312 (N1267, N631, N1159);
MyNand NAND2_313 (N1309, N688, N1205);
MyNand NAND2_314 (N1310, N691, N1207);
MyNand NAND2_315 (N1311, N694, N1209);
MyNand NAND2_316 (N1312, N697, N1211);
MyNand NAND2_317 (N1313, N700, N1213);
MyNand NAND2_318 (N1314, N703, N1215);
MyNand NAND2_319 (N1315, N706, N1220);
MyNand NAND2_320 (N1316, N709, N1223);
MyNand NAND2_321 (N1317, N712, N1225);
MyNand NAND2_322 (N1318, N715, N1228);
MyNot NOT1_323 (N1319, N1158);
MyNand NAND2_324 (N1322, N628, N1230);
MyNand NAND2_325 (N1327, N730, N1238);
MyNand NAND2_326 (N1328, N733, N1241);
MyNot NOT1_327 (N1334, N1162);
MyNand NAND2_328 (N1344, N1267, N1160);
MyNand NAND2_329 (N1345, N1249, N894);
MyNot NOT1_330 (N1346, N1249);
MyNot NOT1_331 (N1348, N1255);
MyNot NOT1_332 (N1349, N1252);
MyNot NOT1_333 (N1350, N1261);
MyNot NOT1_334 (N1351, N1258);
MyNand NAND2_335 (N1352, N1309, N1206);
MyNand NAND2_336 (N1355, N1310, N1208);
MyNand NAND2_337 (N1358, N1311, N1210);
MyNand NAND2_338 (N1361, N1312, N1212);
MyNand NAND2_339 (N1364, N1313, N1214);
MyNand NAND2_340 (N1367, N1314, N1216);
MyNand NAND2_341 (N1370, N1315, N1221);
MyNand NAND2_342 (N1373, N1316, N1224);
MyNand NAND2_343 (N1376, N1317, N1226);
MyNand NAND2_344 (N1379, N1318, N1229);
MyNand NAND2_345 (N1383, N1322, N1231);
MyNot NOT1_346 (N1386, N1232);
MyNand NAND2_347 (N1387, N1232, N990);
MyNot NOT1_348 (N1388, N1235);
MyNand NAND2_349 (N1389, N1235, N993);
MyNand NAND2_350 (N1390, N1327, N1239);
MyNand NAND2_351 (N1393, N1328, N1242);
MyNot NOT1_352 (N1396, N1243);
MyNand NAND2_353 (N1397, N1243, N1004);
MyNot NOT1_354 (N1398, N1246);
MyNand NAND2_355 (N1399, N1246, N1007);
MyNot NOT1_356 (N1409, N1319);
MyNand NAND2_357 (N1412, N649, N1346);
MyNot NOT1_358 (N1413, N1334);
MyBuf BUFF1_359 (N1416, N1264);
MyBuf BUFF1_360 (N1419, N1264);
MyNand NAND2_361 (N1433, N634, N1386);
MyNand NAND2_362 (N1434, N637, N1388);
MyNand NAND2_363 (N1438, N640, N1396);
MyNand NAND2_364 (N1439, N646, N1398);
MyNot NOT1_365 (N1440, N1344);
MyNand NAND2_366 (N1443, N1355, N1148);
MyNot NOT1_367 (N1444, N1355);
MyNand NAND2_368 (N1445, N1352, N1149);
MyNot NOT1_369 (N1446, N1352);
MyNand NAND2_370 (N1447, N1358, N1151);
MyNot NOT1_371 (N1448, N1358);
MyNand NAND2_372 (N1451, N1361, N1152);
MyNot NOT1_373 (N1452, N1361);
MyNand NAND2_374 (N1453, N1367, N1153);
MyNot NOT1_375 (N1454, N1367);
MyNand NAND2_376 (N1455, N1364, N1154);
MyNot NOT1_377 (N1456, N1364);
MyNand NAND2_378 (N1457, N1373, N1156);
MyNot NOT1_379 (N1458, N1373);
MyNand NAND2_380 (N1459, N1379, N1157);
MyNot NOT1_381 (N1460, N1379);
MyNot NOT1_382 (N1461, N1383);
MyNand NAND2_383 (N1462, N1393, N1161);
MyNot NOT1_384 (N1463, N1393);
MyNand NAND2_385 (N1464, N1345, N1412);
MyNot NOT1_386 (N1468, N1370);
MyNand NAND2_387 (N1469, N1370, N1222);
MyNot NOT1_388 (N1470, N1376);
MyNand NAND2_389 (N1471, N1376, N1227);
MyNand NAND2_390 (N1472, N1387, N1433);
MyNot NOT1_391 (N1475, N1390);
MyNand NAND2_392 (N1476, N1390, N1240);
MyNand NAND2_393 (N1478, N1389, N1434);
MyNand NAND2_394 (N1481, N1399, N1439);
MyNand NAND2_395 (N1484, N1397, N1438);
MyNand NAND2_396 (N1487, N939, N1444);
MyNand NAND2_397 (N1488, N935, N1446);
MyNand NAND2_398 (N1489, N943, N1448);
MyNot NOT1_399 (N1490, N1419);
MyNot NOT1_400 (N1491, N1416);
MyNand NAND2_401 (N1492, N947, N1452);
MyNand NAND2_402 (N1493, N955, N1454);
MyNand NAND2_403 (N1494, N951, N1456);
MyNand NAND2_404 (N1495, N969, N1458);
MyNand NAND2_405 (N1496, N977, N1460);
MyNand NAND2_406 (N1498, N998, N1463);
MyNot NOT1_407 (N1499, N1440);
MyNand NAND2_408 (N1500, N965, N1468);
MyNand NAND2_409 (N1501, N973, N1470);
MyNand NAND2_410 (N1504, N994, N1475);
MyNot NOT1_411 (N1510, N1464);
MyNand NAND2_412 (N1513, N1443, N1487);
MyNand NAND2_413 (N1514, N1445, N1488);
MyNand NAND2_414 (N1517, N1447, N1489);
MyNand NAND2_415 (N1520, N1451, N1492);
MyNand NAND2_416 (N1521, N1453, N1493);
MyNand NAND2_417 (N1522, N1455, N1494);
MyNand NAND2_418 (N1526, N1457, N1495);
MyNand NAND2_419 (N1527, N1459, N1496);
MyNot NOT1_420 (N1528, N1472);
MyNand NAND2_421 (N1529, N1462, N1498);
MyNot NOT1_422 (N1530, N1478);
MyNot NOT1_423 (N1531, N1481);
MyNot NOT1_424 (N1532, N1484);
MyNand NAND2_425 (N1534, N1471, N1501);
MyNand NAND2_426 (N1537, N1469, N1500);
MyNand NAND2_427 (N1540, N1476, N1504);
MyNot NOT1_428 (N1546, N1513);
MyNot NOT1_429 (N1554, N1521);
MyNot NOT1_430 (N1557, N1526);
MyNot NOT1_431 (N1561, N1520);
MyNand NAND2_432 (N1567, N1484, N1531);
MyNand NAND2_433 (N1568, N1481, N1532);
MyNot NOT1_434 (N1569, N1510);
MyNot NOT1_435 (N1571, N1527);
MyNot NOT1_436 (N1576, N1529);
MyBuf BUFF1_437 (N1588, N1522);
MyNot NOT1_438 (N1591, N1534);
MyNot NOT1_439 (N1593, N1537);
MyNand NAND2_440 (N1594, N1540, N1530);
MyNot NOT1_441 (N1595, N1540);
MyNand NAND2_442 (N1596, N1567, N1568);
MyBuf BUFF1_443 (N1600, N1517);
MyBuf BUFF1_444 (N1603, N1517);
MyBuf BUFF1_445 (N1606, N1522);
MyBuf BUFF1_446 (N1609, N1522);
MyBuf BUFF1_447 (N1612, N1514);
MyBuf BUFF1_448 (N1615, N1514);
MyBuf BUFF1_449 (N1620, N1557);
MyBuf BUFF1_450 (N1623, N1554);
MyNot NOT1_451 (N1635, N1571);
MyNand NAND2_452 (N1636, N1478, N1595);
MyNand NAND2_453 (N1638, N1576, N1569);
MyNot NOT1_454 (N1639, N1576);
MyBuf BUFF1_455 (N1640, N1561);
MyBuf BUFF1_456 (N1643, N1561);
MyBuf BUFF1_457 (N1647, N1546);
MyBuf BUFF1_458 (N1651, N1546);
MyBuf BUFF1_459 (N1658, N1554);
MyBuf BUFF1_460 (N1661, N1557);
MyBuf BUFF1_461 (N1664, N1557);
MyNand NAND2_462 (N1671, N1596, N893);
MyNot NOT1_463 (N1672, N1596);
MyNot NOT1_464 (N1675, N1600);
MyNot NOT1_465 (N1677, N1603);
MyNand NAND2_466 (N1678, N1606, N1217);
MyNot NOT1_467 (N1679, N1606);
MyNand NAND2_468 (N1680, N1609, N1219);
MyNot NOT1_469 (N1681, N1609);
MyNot NOT1_470 (N1682, N1612);
MyNot NOT1_471 (N1683, N1615);
MyNand NAND2_472 (N1685, N1594, N1636);
MyNand NAND2_473 (N1688, N1510, N1639);
MyBuf BUFF1_474 (N1697, N1588);
MyBuf BUFF1_475 (N1701, N1588);
MyNand NAND2_476 (N1706, N643, N1672);
MyNot NOT1_477 (N1707, N1643);
MyNand NAND2_478 (N1708, N1647, N1675);
MyNot NOT1_479 (N1709, N1647);
MyNand NAND2_480 (N1710, N1651, N1677);
MyNot NOT1_481 (N1711, N1651);
MyNand NAND2_482 (N1712, N1028, N1679);
MyNand NAND2_483 (N1713, N1031, N1681);
MyBuf BUFF1_484 (N1714, N1620);
MyBuf BUFF1_485 (N1717, N1620);
MyNand NAND2_486 (N1720, N1658, N1593);
MyNot NOT1_487 (N1721, N1658);
MyNand NAND2_488 (N1723, N1638, N1688);
MyNot NOT1_489 (N1727, N1661);
MyNot NOT1_490 (N1728, N1640);
MyNot NOT1_491 (N1730, N1664);
MyBuf BUFF1_492 (N1731, N1623);
MyBuf BUFF1_493 (N1734, N1623);
MyNand NAND2_494 (N1740, N1685, N1528);
MyNot NOT1_495 (N1741, N1685);
MyNand NAND2_496 (N1742, N1671, N1706);
MyNand NAND2_497 (N1746, N1600, N1709);
MyNand NAND2_498 (N1747, N1603, N1711);
MyNand NAND2_499 (N1748, N1678, N1712);
MyNand NAND2_500 (N1751, N1680, N1713);
MyNand NAND2_501 (N1759, N1537, N1721);
MyNot NOT1_502 (N1761, N1697);
MyNand NAND2_503 (N1762, N1697, N1727);
MyNot NOT1_504 (N1763, N1701);
MyNand NAND2_505 (N1764, N1701, N1730);
MyNot NOT1_506 (N1768, N1717);
MyNand NAND2_507 (N1769, N1472, N1741);
MyNand NAND2_508 (N1772, N1723, N1413);
MyNot NOT1_509 (N1773, N1723);
MyNand NAND2_510 (N1774, N1708, N1746);
MyNand NAND2_511 (N1777, N1710, N1747);
MyNot NOT1_512 (N1783, N1731);
MyNand NAND2_513 (N1784, N1731, N1682);
MyNot NOT1_514 (N1785, N1714);
MyNot NOT1_515 (N1786, N1734);
MyNand NAND2_516 (N1787, N1734, N1683);
MyNand NAND2_517 (N1788, N1720, N1759);
MyNand NAND2_518 (N1791, N1661, N1761);
MyNand NAND2_519 (N1792, N1664, N1763);
MyNand NAND2_520 (N1795, N1751, N1155);
MyNot NOT1_521 (N1796, N1751);
MyNand NAND2_522 (N1798, N1740, N1769);
MyNand NAND2_523 (N1801, N1334, N1773);
MyNand NAND2_524 (N1802, N1742, N290);
MyNot NOT1_525 (N1807, N1748);
MyNand NAND2_526 (N1808, N1748, N1218);
MyNand NAND2_527 (N1809, N1612, N1783);
MyNand NAND2_528 (N1810, N1615, N1786);
MyNand NAND2_529 (N1812, N1791, N1762);
MyNand NAND2_530 (N1815, N1792, N1764);
MyBuf BUFF1_531 (N1818, N1742);
MyNand NAND2_532 (N1821, N1777, N1490);
MyNot NOT1_533 (N1822, N1777);
MyNand NAND2_534 (N1823, N1774, N1491);
MyNot NOT1_535 (N1824, N1774);
MyNand NAND2_536 (N1825, N962, N1796);
MyNand NAND2_537 (N1826, N1788, N1409);
MyNot NOT1_538 (N1827, N1788);
MyNand NAND2_539 (N1830, N1772, N1801);
MyNand NAND2_540 (N1837, N959, N1807);
MyNand NAND2_541 (N1838, N1809, N1784);
MyNand NAND2_542 (N1841, N1810, N1787);
MyNand NAND2_543 (N1848, N1419, N1822);
MyNand NAND2_544 (N1849, N1416, N1824);
MyNand NAND2_545 (N1850, N1795, N1825);
MyNand NAND2_546 (N1852, N1319, N1827);
MyNand NAND2_547 (N1855, N1815, N1707);
MyNot NOT1_548 (N1856, N1815);
MyNot NOT1_549 (N1857, N1818);
MyNand NAND2_550 (N1858, N1798, N290);
MyNot NOT1_551 (N1864, N1812);
MyNand NAND2_552 (N1865, N1812, N1728);
MyBuf BUFF1_553 (N1866, N1798);
MyBuf BUFF1_554 (N1869, N1802);
MyBuf BUFF1_555 (N1872, N1802);
MyNand NAND2_556 (N1875, N1808, N1837);
MyNand NAND2_557 (N1878, N1821, N1848);
MyNand NAND2_558 (N1879, N1823, N1849);
MyNand NAND2_559 (N1882, N1841, N1768);
MyNot NOT1_560 (N1883, N1841);
MyNand NAND2_561 (N1884, N1826, N1852);
MyNand NAND2_562 (N1885, N1643, N1856);
MyNand NAND2_563 (N1889, N1830, N290);
MyNot NOT1_564 (N1895, N1838);
MyNand NAND2_565 (N1896, N1838, N1785);
MyNand NAND2_566 (N1897, N1640, N1864);
MyNot NOT1_567 (N1898, N1850);
MyBuf BUFF1_568 (N1902, N1830);
MyNot NOT1_569 (N1910, N1878);
MyNand NAND2_570 (N1911, N1717, N1883);
MyNot NOT1_571 (N1912, N1884);
MyNand NAND2_572 (N1913, N1855, N1885);
MyNot NOT1_573 (N1915, N1866);
MyNand NAND2_574 (N1919, N1872, N919);
MyNot NOT1_575 (N1920, N1872);
MyNand NAND2_576 (N1921, N1869, N920);
MyNot NOT1_577 (N1922, N1869);
MyNot NOT1_578 (N1923, N1875);
MyNand NAND2_579 (N1924, N1714, N1895);
MyBuf BUFF1_580 (N1927, N1858);
MyBuf BUFF1_581 (N1930, N1858);
MyNand NAND2_582 (N1933, N1865, N1897);
MyNand NAND2_583 (N1936, N1882, N1911);
MyNot NOT1_584 (N1937, N1898);
MyNot NOT1_585 (N1938, N1902);
MyNand NAND2_586 (N1941, N679, N1920);
MyNand NAND2_587 (N1942, N676, N1922);
MyBuf BUFF1_588 (N1944, N1879);
MyNot NOT1_589 (N1947, N1913);
MyBuf BUFF1_590 (N1950, N1889);
MyBuf BUFF1_591 (N1953, N1889);
MyBuf BUFF1_592 (N1958, N1879);
MyNand NAND2_593 (N1961, N1896, N1924);
MyAnd AND2_594 (N1965, N1910, N601);
MyAnd AND2_595 (N1968, N602, N1912);
MyNand NAND2_596 (N1975, N1930, N917);
MyNot NOT1_597 (N1976, N1930);
MyNand NAND2_598 (N1977, N1927, N918);
MyNot NOT1_599 (N1978, N1927);
MyNand NAND2_600 (N1979, N1919, N1941);
MyNand NAND2_601 (N1980, N1921, N1942);
MyNot NOT1_602 (N1985, N1933);
MyNot NOT1_603 (N1987, N1936);
MyNot NOT1_604 (N1999, N1944);
MyNand NAND2_605 (N2000, N1944, N1937);
MyNot NOT1_606 (N2002, N1947);
MyNand NAND2_607 (N2003, N1947, N1499);
MyNand NAND2_608 (N2004, N1953, N1350);
MyNot NOT1_609 (N2005, N1953);
MyNand NAND2_610 (N2006, N1950, N1351);
MyNot NOT1_611 (N2007, N1950);
MyNand NAND2_612 (N2008, N673, N1976);
MyNand NAND2_613 (N2009, N670, N1978);
MyNot NOT1_614 (N2012, N1979);
MyNot NOT1_615 (N2013, N1958);
MyNand NAND2_616 (N2014, N1958, N1923);
MyNot NOT1_617 (N2015, N1961);
MyNand NAND2_618 (N2016, N1961, N1635);
MyNot NOT1_619 (N2018, N1965);
MyNot NOT1_620 (N2019, N1968);
MyNand NAND2_621 (N2020, N1898, N1999);
MyNot NOT1_622 (N2021, N1987);
MyNand NAND2_623 (N2022, N1987, N1591);
MyNand NAND2_624 (N2023, N1440, N2002);
MyNand NAND2_625 (N2024, N1261, N2005);
MyNand NAND2_626 (N2025, N1258, N2007);
MyNand NAND2_627 (N2026, N1975, N2008);
MyNand NAND2_628 (N2027, N1977, N2009);
MyNot NOT1_629 (N2030, N1980);
MyBuf BUFF1_630 (N2033, N1980);
MyNand NAND2_631 (N2036, N1875, N2013);
MyNand NAND2_632 (N2037, N1571, N2015);
MyNand NAND2_633 (N2038, N2020, N2000);
MyNand NAND2_634 (N2039, N1534, N2021);
MyNand NAND2_635 (N2040, N2023, N2003);
MyNand NAND2_636 (N2041, N2004, N2024);
MyNand NAND2_637 (N2042, N2006, N2025);
MyNot NOT1_638 (N2047, N2026);
MyNand NAND2_639 (N2052, N2036, N2014);
MyNand NAND2_640 (N2055, N2037, N2016);
MyNot NOT1_641 (N2060, N2038);
MyNand NAND2_642 (N2061, N2039, N2022);
MyNand NAND2_643 (N2062, N2040, N290);
MyNot NOT1_644 (N2067, N2041);
MyNot NOT1_645 (N2068, N2027);
MyBuf BUFF1_646 (N2071, N2027);
MyNot NOT1_647 (N2076, N2052);
MyNot NOT1_648 (N2077, N2055);
MyNand NAND2_649 (N2078, N2060, N290);
MyNand NAND2_650 (N2081, N2061, N290);
MyNot NOT1_651 (N2086, N2042);
MyBuf BUFF1_652 (N2089, N2042);
MyAnd AND2_653 (N2104, N2030, N2068);
MyAnd AND2_654 (N2119, N2033, N2068);
MyAnd AND2_655 (N2129, N2030, N2071);
MyAnd AND2_656 (N2143, N2033, N2071);
MyBuf BUFF1_657 (N2148, N2062);
MyBuf BUFF1_658 (N2151, N2062);
MyBuf BUFF1_659 (N2196, N2078);
MyBuf BUFF1_660 (N2199, N2078);
MyBuf BUFF1_661 (N2202, N2081);
MyBuf BUFF1_662 (N2205, N2081);
MyNand NAND2_663 (N2214, N2151, N915);
MyNot NOT1_664 (N2215, N2151);
MyNand NAND2_665 (N2216, N2148, N916);
MyNot NOT1_666 (N2217, N2148);
MyNand NAND2_667 (N2222, N2199, N1348);
MyNot NOT1_668 (N2223, N2199);
MyNand NAND2_669 (N2224, N2196, N1349);
MyNot NOT1_670 (N2225, N2196);
MyNand NAND2_671 (N2226, N2205, N913);
MyNot NOT1_672 (N2227, N2205);
MyNand NAND2_673 (N2228, N2202, N914);
MyNot NOT1_674 (N2229, N2202);
MyNand NAND2_675 (N2230, N667, N2215);
MyNand NAND2_676 (N2231, N664, N2217);
MyNand NAND2_677 (N2232, N1255, N2223);
MyNand NAND2_678 (N2233, N1252, N2225);
MyNand NAND2_679 (N2234, N661, N2227);
MyNand NAND2_680 (N2235, N658, N2229);
MyNand NAND2_681 (N2236, N2214, N2230);
MyNand NAND2_682 (N2237, N2216, N2231);
MyNand NAND2_683 (N2240, N2222, N2232);
MyNand NAND2_684 (N2241, N2224, N2233);
MyNand NAND2_685 (N2244, N2226, N2234);
MyNand NAND2_686 (N2245, N2228, N2235);
MyNot NOT1_687 (N2250, N2236);
MyNot NOT1_688 (N2253, N2240);
MyNot NOT1_689 (N2256, N2244);
MyNot NOT1_690 (N2257, N2237);
MyBuf BUFF1_691 (N2260, N2237);
MyNot NOT1_692 (N2263, N2241);
MyAnd AND2_693 (N2266, N1164, N2241);
MyNot NOT1_694 (N2269, N2245);
MyAnd AND2_695 (N2272, N1168, N2245);
MyNand8 NAND8_696 (N2279, N2067, N2012, N2047, N2250, N899, N2256, N2253, N903);
MyBuf BUFF1_697 (N2286, N2266);
MyBuf BUFF1_698 (N2297, N2266);
MyBuf BUFF1_699 (N2315, N2272);
MyBuf BUFF1_700 (N2326, N2272);
MyAnd AND2_701 (N2340, N2086, N2257);
MyAnd AND2_702 (N2353, N2089, N2257);
MyAnd AND2_703 (N2361, N2086, N2260);
MyAnd AND2_704 (N2375, N2089, N2260);
MyAnd4 AND4_705 (N2384, N338, N2279, N313, N313);
MyAnd AND2_706 (N2385, N1163, N2263);
MyAnd AND2_707 (N2386, N1164, N2263);
MyAnd AND2_708 (N2426, N1167, N2269);
MyAnd AND2_709 (N2427, N1168, N2269);
MyNand5 NAND5_710 (N2537, N2286, N2315, N2361, N2104, N1171);
MyNand5 NAND5_711 (N2540, N2286, N2315, N2340, N2129, N1171);
MyNand5 NAND5_712 (N2543, N2286, N2315, N2340, N2119, N1171);
MyNand5 NAND5_713 (N2546, N2286, N2315, N2353, N2104, N1171);
MyNand5 NAND5_714 (N2549, N2297, N2315, N2375, N2119, N1188);
MyNand5 NAND5_715 (N2552, N2297, N2326, N2361, N2143, N1188);
MyNand5 NAND5_716 (N2555, N2297, N2326, N2375, N2129, N1188);
MyAnd5 AND5_717 (N2558, N2286, N2315, N2361, N2104, N1171);
MyAnd5 AND5_718 (N2561, N2286, N2315, N2340, N2129, N1171);
MyAnd5 AND5_719 (N2564, N2286, N2315, N2340, N2119, N1171);
MyAnd5 AND5_720 (N2567, N2286, N2315, N2353, N2104, N1171);
MyAnd5 AND5_721 (N2570, N2297, N2315, N2375, N2119, N1188);
MyAnd5 AND5_722 (N2573, N2297, N2326, N2361, N2143, N1188);
MyAnd5 AND5_723 (N2576, N2297, N2326, N2375, N2129, N1188);
MyNand5 NAND5_724 (N2594, N2286, N2427, N2361, N2129, N1171);
MyNand5 NAND5_725 (N2597, N2297, N2427, N2361, N2119, N1171);
MyNand5 NAND5_726 (N2600, N2297, N2427, N2375, N2104, N1171);
MyNand5 NAND5_727 (N2603, N2297, N2427, N2340, N2143, N1171);
MyNand5 NAND5_728 (N2606, N2297, N2427, N2353, N2129, N1188);
MyNand5 NAND5_729 (N2611, N2386, N2326, N2361, N2129, N1188);
MyNand5 NAND5_730 (N2614, N2386, N2326, N2361, N2119, N1188);
MyNand5 NAND5_731 (N2617, N2386, N2326, N2375, N2104, N1188);
MyNand5 NAND5_732 (N2620, N2386, N2326, N2353, N2129, N1188);
MyNand5 NAND5_733 (N2627, N2297, N2427, N2340, N2104, N926);
MyNand5 NAND5_734 (N2628, N2386, N2326, N2340, N2104, N926);
MyNand5 NAND5_735 (N2629, N2386, N2427, N2361, N2104, N926);
MyNand5 NAND5_736 (N2630, N2386, N2427, N2340, N2129, N926);
MyNand5 NAND5_737 (N2631, N2386, N2427, N2340, N2119, N926);
MyNand5 NAND5_738 (N2632, N2386, N2427, N2353, N2104, N926);
MyNand5 NAND5_739 (N2633, N2386, N2426, N2340, N2104, N926);
MyNand5 NAND5_740 (N2634, N2385, N2427, N2340, N2104, N926);
MyAnd5 AND5_741 (N2639, N2286, N2427, N2361, N2129, N1171);
MyAnd5 AND5_742 (N2642, N2297, N2427, N2361, N2119, N1171);
MyAnd5 AND5_743 (N2645, N2297, N2427, N2375, N2104, N1171);
MyAnd5 AND5_744 (N2648, N2297, N2427, N2340, N2143, N1171);
MyAnd5 AND5_745 (N2651, N2297, N2427, N2353, N2129, N1188);
MyAnd5 AND5_746 (N2655, N2386, N2326, N2361, N2129, N1188);
MyAnd5 AND5_747 (N2658, N2386, N2326, N2361, N2119, N1188);
MyAnd5 AND5_748 (N2661, N2386, N2326, N2375, N2104, N1188);
MyAnd5 AND5_749 (N2664, N2386, N2326, N2353, N2129, N1188);
MyNand NAND2_750 (N2669, N2558, N534);
MyNot NOT1_751 (N2670, N2558);
MyNand NAND2_752 (N2671, N2561, N535);
MyNot NOT1_753 (N2672, N2561);
MyNand NAND2_754 (N2673, N2564, N536);
MyNot NOT1_755 (N2674, N2564);
MyNand NAND2_756 (N2675, N2567, N537);
MyNot NOT1_757 (N2676, N2567);
MyNand NAND2_758 (N2682, N2570, N543);
MyNot NOT1_759 (N2683, N2570);
MyNand NAND2_760 (N2688, N2573, N548);
MyNot NOT1_761 (N2689, N2573);
MyNand NAND2_762 (N2690, N2576, N549);
MyNot NOT1_763 (N2691, N2576);
MyAnd8 AND8_764 (N2710, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634);
MyNand NAND2_765 (N2720, N343, N2670);
MyNand NAND2_766 (N2721, N346, N2672);
MyNand NAND2_767 (N2722, N349, N2674);
MyNand NAND2_768 (N2723, N352, N2676);
MyNand NAND2_769 (N2724, N2639, N538);
MyNot NOT1_770 (N2725, N2639);
MyNand NAND2_771 (N2726, N2642, N539);
MyNot NOT1_772 (N2727, N2642);
MyNand NAND2_773 (N2728, N2645, N540);
MyNot NOT1_774 (N2729, N2645);
MyNand NAND2_775 (N2730, N2648, N541);
MyNot NOT1_776 (N2731, N2648);
MyNand NAND2_777 (N2732, N2651, N542);
MyNot NOT1_778 (N2733, N2651);
MyNand NAND2_779 (N2734, N370, N2683);
MyNand NAND2_780 (N2735, N2655, N544);
MyNot NOT1_781 (N2736, N2655);
MyNand NAND2_782 (N2737, N2658, N545);
MyNot NOT1_783 (N2738, N2658);
MyNand NAND2_784 (N2739, N2661, N546);
MyNot NOT1_785 (N2740, N2661);
MyNand NAND2_786 (N2741, N2664, N547);
MyNot NOT1_787 (N2742, N2664);
MyNand NAND2_788 (N2743, N385, N2689);
MyNand NAND2_789 (N2744, N388, N2691);
MyNand8 NAND8_790 (N2745, N2537, N2540, N2543, N2546, N2594, N2597, N2600, N2603);
MyNand8 NAND8_791 (N2746, N2606, N2549, N2611, N2614, N2617, N2620, N2552, N2555);
MyAnd8 AND8_792 (N2747, N2537, N2540, N2543, N2546, N2594, N2597, N2600, N2603);
MyAnd8 AND8_793 (N2750, N2606, N2549, N2611, N2614, N2617, N2620, N2552, N2555);
MyNand NAND2_794 (N2753, N2669, N2720);
MyNand NAND2_795 (N2754, N2671, N2721);
MyNand NAND2_796 (N2755, N2673, N2722);
MyNand NAND2_797 (N2756, N2675, N2723);
MyNand NAND2_798 (N2757, N355, N2725);
MyNand NAND2_799 (N2758, N358, N2727);
MyNand NAND2_800 (N2759, N361, N2729);
MyNand NAND2_801 (N2760, N364, N2731);
MyNand NAND2_802 (N2761, N367, N2733);
MyNand NAND2_803 (N2762, N2682, N2734);
MyNand NAND2_804 (N2763, N373, N2736);
MyNand NAND2_805 (N2764, N376, N2738);
MyNand NAND2_806 (N2765, N379, N2740);
MyNand NAND2_807 (N2766, N382, N2742);
MyNand NAND2_808 (N2767, N2688, N2743);
MyNand NAND2_809 (N2768, N2690, N2744);
MyAnd AND2_810 (N2773, N2745, N275);
MyAnd AND2_811 (N2776, N2746, N276);
MyNand NAND2_812 (N2779, N2724, N2757);
MyNand NAND2_813 (N2780, N2726, N2758);
MyNand NAND2_814 (N2781, N2728, N2759);
MyNand NAND2_815 (N2782, N2730, N2760);
MyNand NAND2_816 (N2783, N2732, N2761);
MyNand NAND2_817 (N2784, N2735, N2763);
MyNand NAND2_818 (N2785, N2737, N2764);
MyNand NAND2_819 (N2786, N2739, N2765);
MyNand NAND2_820 (N2787, N2741, N2766);
MyAnd3 AND3_821 (N2788, N2747, N2750, N2710);
MyNand NAND2_822 (N2789, N2747, N2750);
MyAnd4 AND4_823 (N2800, N338, N2279, N99, N2788);
MyNand NAND2_824 (N2807, N2773, N2018);
MyNot NOT1_825 (N2808, N2773);
MyNand NAND2_826 (N2809, N2776, N2019);
MyNot NOT1_827 (N2810, N2776);
MyNor NOR2_828 (N2811, N2384, N2800);
MyAnd3 AND3_829 (N2812, N897, N283, N2789);
MyAnd3 AND3_830 (N2815, N76, N283, N2789);
MyAnd3 AND3_831 (N2818, N82, N283, N2789);
MyAnd3 AND3_832 (N2821, N85, N283, N2789);
MyAnd3 AND3_833 (N2824, N898, N283, N2789);
MyNand NAND2_834 (N2827, N1965, N2808);
MyNand NAND2_835 (N2828, N1968, N2810);
MyAnd3 AND3_836 (N2829, N79, N283, N2789);
MyNand NAND2_837 (N2843, N2807, N2827);
MyNand NAND2_838 (N2846, N2809, N2828);
MyNand NAND2_839 (N2850, N2812, N2076);
MyNand NAND2_840 (N2851, N2815, N2077);
MyNand NAND2_841 (N2852, N2818, N1915);
MyNand NAND2_842 (N2853, N2821, N1857);
MyNand NAND2_843 (N2854, N2824, N1938);
MyNot NOT1_844 (N2857, N2812);
MyNot NOT1_845 (N2858, N2815);
MyNot NOT1_846 (N2859, N2818);
MyNot NOT1_847 (N2860, N2821);
MyNot NOT1_848 (N2861, N2824);
MyNot NOT1_849 (N2862, N2829);
MyNand NAND2_850 (N2863, N2829, N1985);
MyNand NAND2_851 (N2866, N2052, N2857);
MyNand NAND2_852 (N2867, N2055, N2858);
MyNand NAND2_853 (N2868, N1866, N2859);
MyNand NAND2_854 (N2869, N1818, N2860);
MyNand NAND2_855 (N2870, N1902, N2861);
MyNand NAND2_856 (N2871, N2843, N886);
MyNot NOT1_857 (N2872, N2843);
MyNand NAND2_858 (N2873, N2846, N887);
MyNot NOT1_859 (N2874, N2846);
MyNand NAND2_860 (N2875, N1933, N2862);
MyNand NAND2_861 (N2876, N2866, N2850);
MyNand NAND2_862 (N2877, N2867, N2851);
MyNand NAND2_863 (N2878, N2868, N2852);
MyNand NAND2_864 (N2879, N2869, N2853);
MyNand NAND2_865 (N2880, N2870, N2854);
MyNand NAND2_866 (N2881, N682, N2872);
MyNand NAND2_867 (N2882, N685, N2874);
MyNand NAND2_868 (N2883, N2875, N2863);
MyAnd AND2_869 (N2886, N2876, N550);
MyAnd AND2_870 (N2887, N551, N2877);
MyAnd AND2_871 (N2888, N553, N2878);
MyAnd AND2_872 (N2889, N2879, N554);
MyAnd AND2_873 (N2890, N555, N2880);
MyNand NAND2_874 (N2891, N2871, N2881);
MyNand NAND2_875 (N2892, N2873, N2882);
MyNand NAND2_876 (N2895, N2883, N1461);
MyNot NOT1_877 (N2896, N2883);
MyNand NAND2_878 (N2897, N1383, N2896);
MyNand NAND2_879 (N2898, N2895, N2897);
MyAnd AND2_880 (N2899, N2898, N552);

endmodule
